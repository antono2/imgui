@[translated]
module implot

#flag -I @VMODROOT/include

#include <time.h>

#include <cimplot.h>

#flag -DIMGUI_USE_WCHAR32

pub struct InputMap {
	pan           ImGuiMouseButton
	panMod        int
	fit           ImGuiMouseButton
	select        ImGuiMouseButton
	selectCancel  ImGuiMouseButton
	selectMod     int
	selectHorzMod int
	selectVertMod int
	menu          ImGuiMouseButton
	overrideMod   int
	zoomMod       int
	zoomRate      f32
}

pub type C.tm = voidptr

pub type C.time_t = voidptr

// This file is automatically generated by int(generator.lua) from https://int(github.com)/cimgui/cimgui
// based on int(imgui.h) file version "1.91.9b" 19191 from Dear ImGui https://int(github.com)/ocornut/imgui
// with int(imgui_internal.h) api
// with int(imgui_freetype.h) api
// docking branch
// typedef unsigned long long ImU64;
struct ImVector_const_charPtr {
	size     int
	capacity int
	data     &&u8
}

type ImGuiID = u32
type ImS8 = i8
type ImU8 = u8
type ImS16 = i16
type ImU16 = u16
type ImS32 = int
type ImU32 = u32
type ImS64 = i64
type ImU64 = i64
type ImGuiCol = int
type ImGuiCond = int
type ImGuiDataType = int
type ImGuiMouseButton = int
type ImGuiMouseCursor = int
type ImGuiStyleVar = int
type ImGuiTableBgTarget = int
type ImDrawFlags = int
type ImDrawListFlags = int
type ImFontAtlasFlags = int
type ImGuiBackendFlags = int
type ImGuiButtonFlags = int
type ImGuiChildFlags = int
type ImGuiColorEditFlags = int
type ImGuiConfigFlags = int
type ImGuiComboFlags = int
type ImGuiDockNodeFlags = int
type ImGuiDragDropFlags = int
type ImGuiFocusedFlags = int
type ImGuiHoveredFlags = int
type ImGuiInputFlags = int
type ImGuiInputTextFlags = int
type ImGuiItemFlags = int
type ImGuiKeyChord = int
type ImGuiPopupFlags = int
type ImGuiMultiSelectFlags = int
type ImGuiSelectableFlags = int
type ImGuiSliderFlags = int
type ImGuiTabBarFlags = int
type ImGuiTabItemFlags = int
type ImGuiTableFlags = int
type ImGuiTableColumnFlags = int
type ImGuiTableRowFlags = int
type ImGuiTreeNodeFlags = int
type ImGuiViewportFlags = int
type ImGuiWindowFlags = int
type ImWchar32 = u32
type ImWchar16 = u16
type ImGuiSelectionUserData = i64
type ImGuiMemAllocFunc = fn (usize, voidptr) voidptr

type ImGuiMemFreeFunc = fn (voidptr, voidptr)

struct ImVec2 {
	x f32
	y f32
}

struct ImTextureID {
	x f32
	y f32
	z f32
	w f32
}

enum ImGuiWindowFlags_ {
	none                        = 0
	no_title_bar                = 1 << 0
	no_resize                   = 1 << 1
	no_move                     = 1 << 2
	no_scrollbar                = 1 << 3
	no_scroll_with_mouse        = 1 << 4
	no_collapse                 = 1 << 5
	always_auto_resize          = 1 << 6
	no_background               = 1 << 7
	no_saved_settings           = 1 << 8
	no_mouse_inputs             = 1 << 9
	menu_bar                    = 1 << 10
	horizontal_scrollbar        = 1 << 11
	no_focus_on_appearing       = 1 << 12
	no_bring_to_front_on_focus  = 1 << 13
	always_vertical_scrollbar   = 1 << 14
	always_horizontal_scrollbar = 1 << 15
	no_nav_inputs               = 1 << 16
	no_nav_focus                = 1 << 17
	unsaved_document            = 1 << 18
	no_docking                  = 1 << 19
	no_nav                      = 1 << 16 | 1 << 17
	no_decoration               = 1 << 0 | 1 << 1 | 1 << 3 | 1 << 5
	no_inputs                   = 1 << 9 | 1 << 16 | 1 << 17
	dock_node_host              = 1 << 23
	child_window                = 1 << 24
	tooltip                     = 1 << 25
	popup                       = 1 << 26
	modal                       = 1 << 27
	child_menu                  = 1 << 28
}

enum ImGuiChildFlags_ {
	none                      = 0
	borders                   = 1 << 0
	always_use_window_padding = 1 << 1
	resize_x                  = 1 << 2
	resize_y                  = 1 << 3
	auto_resize_x             = 1 << 4
	auto_resize_y             = 1 << 5
	always_auto_resize        = 1 << 6
	frame_style               = 1 << 7
	nav_flattened             = 1 << 8
}

enum ImGuiItemFlags_ {
	none                 = 0
	no_tab_stop          = 1 << 0
	no_nav               = 1 << 1
	no_nav_default_focus = 1 << 2
	button_repeat        = 1 << 3
	auto_close_popups    = 1 << 4
	allow_duplicate_id   = 1 << 5
}

enum ImGuiInputTextFlags_ {
	none                    = 0
	chars_decimal           = 1 << 0
	chars_hexadecimal       = 1 << 1
	chars_scientific        = 1 << 2
	chars_uppercase         = 1 << 3
	chars_no_blank          = 1 << 4
	allow_tab_input         = 1 << 5
	enter_returns_true      = 1 << 6
	escape_clears_all       = 1 << 7
	ctrl_enter_for_new_line = 1 << 8
	read_only               = 1 << 9
	password                = 1 << 10
	always_overwrite        = 1 << 11
	auto_select_all         = 1 << 12
	parse_empty_ref_val     = 1 << 13
	display_empty_ref_val   = 1 << 14
	no_horizontal_scroll    = 1 << 15
	no_undo_redo            = 1 << 16
	elide_left              = 1 << 17
	callback_completion     = 1 << 18
	callback_history        = 1 << 19
	callback_always         = 1 << 20
	callback_char_filter    = 1 << 21
	callback_resize         = 1 << 22
	callback_edit           = 1 << 23
}

enum ImGuiTreeNodeFlags_ {
	none                     = 0
	selected                 = 1 << 0
	framed                   = 1 << 1
	allow_overlap            = 1 << 2
	no_tree_push_on_open     = 1 << 3
	no_auto_open_on_log      = 1 << 4
	default_open             = 1 << 5
	open_on_double_click     = 1 << 6
	open_on_arrow            = 1 << 7
	leaf                     = 1 << 8
	bullet                   = 1 << 9
	frame_padding            = 1 << 10
	span_avail_width         = 1 << 11
	span_full_width          = 1 << 12
	span_label_width         = 1 << 13
	span_all_columns         = 1 << 14
	label_span_all_columns   = 1 << 15
	nav_left_jumps_back_here = 1 << 17
	collapsing_header        = 1 << 1 | 1 << 3 | 1 << 4
}

enum ImGuiPopupFlags_ {
	none                        = 0
	mouse_button_left           = 0
	mouse_button_right          = 1
	mouse_button_middle         = 2
	mouse_button_mask_          = 31
	mouse_button_default_       = 1
	no_reopen                   = 1 << 5
	no_open_over_existing_popup = 1 << 7
	no_open_over_items          = 1 << 8
	any_popup_id                = 1 << 10
	any_popup_level             = 1 << 11
	any_popup                   = 1 << 10 | 1 << 11
}

enum ImGuiSelectableFlags_ {
	none                 = 0
	no_auto_close_popups = 1 << 0
	span_all_columns     = 1 << 1
	allow_double_click   = 1 << 2
	disabled             = 1 << 3
	allow_overlap        = 1 << 4
	highlight            = 1 << 5
}

enum ImGuiComboFlags_ {
	none              = 0
	popup_align_left  = 1 << 0
	height_small      = 1 << 1
	height_regular    = 1 << 2
	height_large      = 1 << 3
	height_largest    = 1 << 4
	no_arrow_button   = 1 << 5
	no_preview        = 1 << 6
	width_fit_preview = 1 << 7
	height_mask_      = 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4
}

enum ImGuiTabBarFlags_ {
	none                              = 0
	reorderable                       = 1 << 0
	auto_select_new_tabs              = 1 << 1
	tab_list_popup_button             = 1 << 2
	no_close_with_middle_mouse_button = 1 << 3
	no_tab_list_scrolling_buttons     = 1 << 4
	no_tooltip                        = 1 << 5
	draw_selected_overline            = 1 << 6
	fitting_policy_resize_down        = 1 << 7
	fitting_policy_scroll             = 1 << 8
	fitting_policy_mask_              = 1 << 7 | 1 << 8
	fitting_policy_default_           = 1 << 7
}

enum ImGuiTabItemFlags_ {
	none                              = 0
	unsaved_document                  = 1 << 0
	set_selected                      = 1 << 1
	no_close_with_middle_mouse_button = 1 << 2
	no_push_id                        = 1 << 3
	no_tooltip                        = 1 << 4
	no_reorder                        = 1 << 5
	leading                           = 1 << 6
	trailing                          = 1 << 7
	no_assumed_closure                = 1 << 8
}

enum ImGuiFocusedFlags_ {
	none                   = 0
	child_windows          = 1 << 0
	root_window            = 1 << 1
	any_window             = 1 << 2
	no_popup_hierarchy     = 1 << 3
	dock_hierarchy         = 1 << 4
	root_and_child_windows = 1 << 1 | 1 << 0
}

enum ImGuiHoveredFlags_ {
	none                              = 0
	child_windows                     = 1 << 0
	root_window                       = 1 << 1
	any_window                        = 1 << 2
	no_popup_hierarchy                = 1 << 3
	dock_hierarchy                    = 1 << 4
	allow_when_blocked_by_popup       = 1 << 5
	allow_when_blocked_by_active_item = 1 << 7
	allow_when_overlapped_by_item     = 1 << 8
	allow_when_overlapped_by_window   = 1 << 9
	allow_when_disabled               = 1 << 10
	no_nav_override                   = 1 << 11
	allow_when_overlapped             = 1 << 8 | 1 << 9
	rect_only                         = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9
	root_and_child_windows            = 1 << 1 | 1 << 0
	for_tooltip                       = 1 << 12
	stationary                        = 1 << 13
	delay_none                        = 1 << 14
	delay_short                       = 1 << 15
	delay_normal                      = 1 << 16
	no_shared_delay                   = 1 << 17
}

enum ImGuiDockNodeFlags_ {
	none                         = 0
	keep_alive_only              = 1 << 0
	no_docking_over_central_node = 1 << 2
	passthru_central_node        = 1 << 3
	no_docking_split             = 1 << 4
	no_resize                    = 1 << 5
	auto_hide_tab_bar            = 1 << 6
	no_undocking                 = 1 << 7
}

enum ImGuiDragDropFlags_ {
	none                          = 0
	source_no_preview_tooltip     = 1 << 0
	source_no_disable_hover       = 1 << 1
	source_no_hold_to_open_others = 1 << 2
	source_allow_null_id          = 1 << 3
	source_extern                 = 1 << 4
	payload_auto_expire           = 1 << 5
	payload_no_cross_context      = 1 << 6
	payload_no_cross_process      = 1 << 7
	accept_before_delivery        = 1 << 10
	accept_no_draw_default_rect   = 1 << 11
	accept_no_preview_tooltip     = 1 << 12
	accept_peek_only              = 1 << 10 | 1 << 11
}

enum ImGuiDataType_ {
	s8
	u8
	s16
	u16
	s32
	u32
	s64
	u64
	float
	double
	bool
	string
	count
}

enum ImGuiDir {
	none  = -1
	left  = 0
	right = 1
	up    = 2
	down  = 3
	count = 4
}

enum ImGuiSortDirection {
	none       = 0
	ascending  = 1
	descending = 2
}

enum ImGuiKey {
	none                   = 0
	named_begin            = 512
	tab                    = 512
	left_arrow             = 513
	right_arrow            = 514
	up_arrow               = 515
	down_arrow             = 516
	page_up                = 517
	page_down              = 518
	home                   = 519
	end                    = 520
	insert                 = 521
	delete                 = 522
	backspace              = 523
	space                  = 524
	enter                  = 525
	escape                 = 526
	left_ctrl              = 527
	left_shift             = 528
	left_alt               = 529
	left_super             = 530
	right_ctrl             = 531
	right_shift            = 532
	right_alt              = 533
	right_super            = 534
	menu                   = 535
	_0                     = 536
	_1                     = 537
	_2                     = 538
	_3                     = 539
	_4                     = 540
	_5                     = 541
	_6                     = 542
	_7                     = 543
	_8                     = 544
	_9                     = 545
	a                      = 546
	b                      = 547
	c                      = 548
	d                      = 549
	e                      = 550
	f                      = 551
	g                      = 552
	h                      = 553
	i                      = 554
	j                      = 555
	k                      = 556
	l                      = 557
	m                      = 558
	n                      = 559
	o                      = 560
	p                      = 561
	q                      = 562
	r                      = 563
	s                      = 564
	t                      = 565
	u                      = 566
	v                      = 567
	w                      = 568
	x                      = 569
	y                      = 570
	z                      = 571
	f1                     = 572
	f2                     = 573
	f3                     = 574
	f4                     = 575
	f5                     = 576
	f6                     = 577
	f7                     = 578
	f8                     = 579
	f9                     = 580
	f10                    = 581
	f11                    = 582
	f12                    = 583
	f13                    = 584
	f14                    = 585
	f15                    = 586
	f16                    = 587
	f17                    = 588
	f18                    = 589
	f19                    = 590
	f20                    = 591
	f21                    = 592
	f22                    = 593
	f23                    = 594
	f24                    = 595
	apostrophe             = 596
	comma                  = 597
	minus                  = 598
	period                 = 599
	slash                  = 600
	semicolon              = 601
	equal                  = 602
	left_bracket           = 603
	backslash              = 604
	right_bracket          = 605
	grave_accent           = 606
	caps_lock              = 607
	scroll_lock            = 608
	num_lock               = 609
	print_screen           = 610
	pause                  = 611
	pad0                   = 612
	pad1                   = 613
	pad2                   = 614
	pad3                   = 615
	pad4                   = 616
	pad5                   = 617
	pad6                   = 618
	pad7                   = 619
	pad8                   = 620
	pad9                   = 621
	pad_decimal            = 622
	pad_divide             = 623
	pad_multiply           = 624
	pad_subtract           = 625
	pad_add                = 626
	pad_enter              = 627
	pad_equal              = 628
	app_back               = 629
	app_forward            = 630
	oem102                 = 631
	gamepad_start          = 632
	gamepad_back           = 633
	gamepad_face_left      = 634
	gamepad_face_right     = 635
	gamepad_face_up        = 636
	gamepad_face_down      = 637
	gamepad_dpad_left      = 638
	gamepad_dpad_right     = 639
	gamepad_dpad_up        = 640
	gamepad_dpad_down      = 641
	gamepad_l1             = 642
	gamepad_r1             = 643
	gamepad_l2             = 644
	gamepad_r2             = 645
	gamepad_l3             = 646
	gamepad_r3             = 647
	gamepad_ls_tick_left   = 648
	gamepad_ls_tick_right  = 649
	gamepad_ls_tick_up     = 650
	gamepad_ls_tick_down   = 651
	gamepad_rs_tick_left   = 652
	gamepad_rs_tick_right  = 653
	gamepad_rs_tick_up     = 654
	gamepad_rs_tick_down   = 655
	mouse_left             = 656
	mouse_right            = 657
	mouse_middle           = 658
	mouse_x1               = 659
	mouse_x2               = 660
	mouse_wheel_x          = 661
	mouse_wheel_y          = 662
	reserved_for_mod_ctrl  = 663
	reserved_for_mod_shift = 664
	reserved_for_mod_alt   = 665
	reserved_for_mod_super = 666
	named_end              = 667
	mod_none               = 0
	mod_ctrl               = 1 << 12
	mod_shift              = 1 << 13
	mod_alt                = 1 << 14
	mod_super              = 1 << 15
	mod_mask_              = 61440
	named_count            = 667 - 512
}

enum ImGuiInputFlags_ {
	none                    = 0
	repeat                  = 1 << 0
	route_active            = 1 << 10
	route_focused           = 1 << 11
	route_global            = 1 << 12
	route_always            = 1 << 13
	route_over_focused      = 1 << 14
	route_over_active       = 1 << 15
	route_unless_bg_focused = 1 << 16
	route_from_root_window  = 1 << 17
	tooltip                 = 1 << 18
}

enum ImGuiConfigFlags_ {
	none                       = 0
	nav_enable_keyboard        = 1 << 0
	nav_enable_gamepad         = 1 << 1
	no_mouse                   = 1 << 4
	no_mouse_cursor_change     = 1 << 5
	no_keyboard                = 1 << 6
	docking_enable             = 1 << 7
	viewports_enable           = 1 << 10
	dpi_enable_scale_viewports = 1 << 14
	dpi_enable_scale_fonts     = 1 << 15
	is_srgb                    = 1 << 20
	is_touch_screen            = 1 << 21
}

enum ImGuiBackendFlags_ {
	none                       = 0
	has_gamepad                = 1 << 0
	has_mouse_cursors          = 1 << 1
	has_set_mouse_pos          = 1 << 2
	renderer_has_vtx_offset    = 1 << 3
	platform_has_viewports     = 1 << 10
	has_mouse_hovered_viewport = 1 << 11
	renderer_has_viewports     = 1 << 12
}

enum ImGuiCol_ {
	text
	text_disabled
	window_bg
	child_bg
	popup_bg
	border
	border_shadow
	frame_bg
	frame_bg_hovered
	frame_bg_active
	title_bg
	title_bg_active
	title_bg_collapsed
	menu_bar_bg
	scrollbar_bg
	scrollbar_grab
	scrollbar_grab_hovered
	scrollbar_grab_active
	check_mark
	slider_grab
	slider_grab_active
	button
	button_hovered
	button_active
	header
	header_hovered
	header_active
	separator
	separator_hovered
	separator_active
	resize_grip
	resize_grip_hovered
	resize_grip_active
	tab_hovered
	tab
	tab_selected
	tab_selected_overline
	tab_dimmed
	tab_dimmed_selected
	tab_dimmed_selected_overline
	docking_preview
	docking_empty_bg
	plot_lines
	plot_lines_hovered
	plot_histogram
	plot_histogram_hovered
	table_header_bg
	table_border_strong
	table_border_light
	table_row_bg
	table_row_bg_alt
	text_link
	text_selected_bg
	drag_drop_target
	nav_cursor
	nav_windowing_highlight
	nav_windowing_dim_bg
	modal_window_dim_bg
	count
}

enum ImGuiStyleVar_ {
	alpha
	disabled_alpha
	window_padding
	window_rounding
	window_border_size
	window_min_size
	window_title_align
	child_rounding
	child_border_size
	popup_rounding
	popup_border_size
	frame_padding
	frame_rounding
	frame_border_size
	item_spacing
	item_inner_spacing
	indent_spacing
	cell_padding
	scrollbar_size
	scrollbar_rounding
	grab_min_size
	grab_rounding
	image_border_size
	tab_rounding
	tab_border_size
	tab_bar_border_size
	tab_bar_overline_size
	table_angled_headers_angle
	table_angled_headers_text_align
	button_text_align
	selectable_text_align
	separator_text_border_size
	separator_text_align
	separator_text_padding
	docking_separator_size
	count
}

enum ImGuiButtonFlags_ {
	none                = 0
	mouse_button_left   = 1 << 0
	mouse_button_right  = 1 << 1
	mouse_button_middle = 1 << 2
	mouse_button_mask_  = 1 << 0 | 1 << 1 | 1 << 2
	enable_nav          = 1 << 3
}

enum ImGuiColorEditFlags_ {
	none               = 0
	no_alpha           = 1 << 1
	no_picker          = 1 << 2
	no_options         = 1 << 3
	no_small_preview   = 1 << 4
	no_inputs          = 1 << 5
	no_tooltip         = 1 << 6
	no_label           = 1 << 7
	no_side_preview    = 1 << 8
	no_drag_drop       = 1 << 9
	no_border          = 1 << 10
	alpha_opaque       = 1 << 11
	alpha_no_bg        = 1 << 12
	alpha_preview_half = 1 << 13
	alpha_bar          = 1 << 16
	hdr                = 1 << 19
	display_rgb        = 1 << 20
	display_hsv        = 1 << 21
	display_hex        = 1 << 22
	uint8              = 1 << 23
	float              = 1 << 24
	picker_hue_bar     = 1 << 25
	picker_hue_wheel   = 1 << 26
	input_rgb          = 1 << 27
	input_hsv          = 1 << 28
	default_options_   = 1 << 23 | 1 << 20 | 1 << 27 | 1 << 25
	alpha_mask_        = 1 << 1 | 1 << 11 | 1 << 12 | 1 << 13
	display_mask_      = 1 << 20 | 1 << 21 | 1 << 22
	data_type_mask_    = 1 << 23 | 1 << 24
	picker_mask_       = 1 << 26 | 1 << 25
	input_mask_        = 1 << 27 | 1 << 28
}

enum ImGuiSliderFlags_ {
	none               = 0
	logarithmic        = 1 << 5
	no_round_to_format = 1 << 6
	no_input           = 1 << 7
	wrap_around        = 1 << 8
	clamp_on_input     = 1 << 9
	clamp_zero_range   = 1 << 10
	no_speed_tweaks    = 1 << 11
	always_clamp       = 1 << 9 | 1 << 10
	invalid_mask_      = 1879048207
}

enum ImGuiMouseButton_ {
	left   = 0
	right  = 1
	middle = 2
	count  = 5
}

enum ImGuiMouseCursor_ {
	none  = -1
	arrow = 0
	text_input
	resize_all
	resize_ns
	resize_ew
	resize_nesw
	resize_nwse
	hand
	wait
	progress
	not_allowed
	count
}

enum ImGuiMouseSource {
	mouse        = 0
	touch_screen = 1
	pen          = 2
	count        = 3
}

enum ImGuiCond_ {
	none           = 0
	always         = 1 << 0
	once           = 1 << 1
	first_use_ever = 1 << 2
	appearing      = 1 << 3
}

enum ImGuiTableFlags_ {
	none                            = 0
	resizable                       = 1 << 0
	reorderable                     = 1 << 1
	hideable                        = 1 << 2
	sortable                        = 1 << 3
	no_saved_settings               = 1 << 4
	context_menu_in_body            = 1 << 5
	row_bg                          = 1 << 6
	borders_inner_h                 = 1 << 7
	borders_outer_h                 = 1 << 8
	borders_inner_v                 = 1 << 9
	borders_outer_v                 = 1 << 10
	borders_h                       = 1 << 7 | 1 << 8
	borders_v                       = 1 << 9 | 1 << 10
	borders_inner                   = 1 << 9 | 1 << 7
	borders_outer                   = 1 << 10 | 1 << 8
	borders                         = 1 << 9 | 1 << 7 | 1 << 10 | 1 << 8
	no_borders_in_body              = 1 << 11
	no_borders_in_body_until_resize = 1 << 12
	sizing_fixed_fit                = 1 << 13
	sizing_fixed_same               = 2 << 13
	sizing_stretch_prop             = 3 << 13
	sizing_stretch_same             = 4 << 13
	no_host_extend_x                = 1 << 16
	no_host_extend_y                = 1 << 17
	no_keep_columns_visible         = 1 << 18
	precise_widths                  = 1 << 19
	no_clip                         = 1 << 20
	pad_outer_x                     = 1 << 21
	no_pad_outer_x                  = 1 << 22
	no_pad_inner_x                  = 1 << 23
	scroll_x                        = 1 << 24
	scroll_y                        = 1 << 25
	sort_multi                      = 1 << 26
	sort_tristate                   = 1 << 27
	highlight_hovered_column        = 1 << 28
	sizing_mask_                    = 1 << 13 | 2 << 13 | 3 << 13 | 4 << 13
}

enum ImGuiTableColumnFlags_ {
	none                   = 0
	disabled               = 1 << 0
	default_hide           = 1 << 1
	default_sort           = 1 << 2
	width_stretch          = 1 << 3
	width_fixed            = 1 << 4
	no_resize              = 1 << 5
	no_reorder             = 1 << 6
	no_hide                = 1 << 7
	no_clip                = 1 << 8
	no_sort                = 1 << 9
	no_sort_ascending      = 1 << 10
	no_sort_descending     = 1 << 11
	no_header_label        = 1 << 12
	no_header_width        = 1 << 13
	prefer_sort_ascending  = 1 << 14
	prefer_sort_descending = 1 << 15
	indent_enable          = 1 << 16
	indent_disable         = 1 << 17
	angled_header          = 1 << 18
	is_enabled             = 1 << 24
	is_visible             = 1 << 25
	is_sorted              = 1 << 26
	is_hovered             = 1 << 27
	width_mask_            = 1 << 3 | 1 << 4
	indent_mask_           = 1 << 16 | 1 << 17
	status_mask_           = 1 << 24 | 1 << 25 | 1 << 26 | 1 << 27
	no_direct_resize_      = 1 << 30
}

enum ImGuiTableRowFlags_ {
	none    = 0
	headers = 1 << 0
}

enum ImGuiTableBgTarget_ {
	none    = 0
	row_bg0 = 1
	row_bg1 = 2
	cell_bg = 3
}

struct ImGuiTableSortSpecs {
	specs      &ImGuiTableColumnSortSpecs
	specsCount int
	specsDirty bool
}

struct ImGuiTableColumnSortSpecs {
	columnUserID  ImGuiID
	columnIndex   ImS16
	sortOrder     ImS16
	sortDirection ImGuiSortDirection
}

struct ImGuiStyle {
	alpha                            f32
	disabledAlpha                    f32
	windowPadding                    ImVec2
	windowRounding                   f32
	windowBorderSize                 f32
	windowBorderHoverPadding         f32
	windowMinSize                    ImVec2
	windowTitleAlign                 ImVec2
	windowMenuButtonPosition         ImGuiDir
	childRounding                    f32
	childBorderSize                  f32
	popupRounding                    f32
	popupBorderSize                  f32
	framePadding                     ImVec2
	frameRounding                    f32
	frameBorderSize                  f32
	itemSpacing                      ImVec2
	itemInnerSpacing                 ImVec2
	cellPadding                      ImVec2
	touchExtraPadding                ImVec2
	indentSpacing                    f32
	columnsMinSpacing                f32
	scrollbarSize                    f32
	scrollbarRounding                f32
	grabMinSize                      f32
	grabRounding                     f32
	logSliderDeadzone                f32
	imageBorderSize                  f32
	tabRounding                      f32
	tabBorderSize                    f32
	tabCloseButtonMinWidthSelected   f32
	tabCloseButtonMinWidthUnselected f32
	tabBarBorderSize                 f32
	tabBarOverlineSize               f32
	tableAngledHeadersAngle          f32
	tableAngledHeadersTextAlign      ImVec2
	colorButtonPosition              ImGuiDir
	buttonTextAlign                  ImVec2
	selectableTextAlign              ImVec2
	separatorTextBorderSize          f32
	separatorTextAlign               ImVec2
	separatorTextPadding             ImVec2
	displayWindowPadding             ImVec2
	displaySafeAreaPadding           ImVec2
	dockingSeparatorSize             f32
	mouseCursorScale                 f32
	antiAliasedLines                 bool
	antiAliasedLinesUseTex           bool
	antiAliasedFill                  bool
	curveTessellationTol             f32
	circleTessellationMaxError       f32
	colors                           [58]C.ImVec4
	hoverStationaryDelay             f32
	hoverDelayShort                  f32
	hoverDelayNormal                 f32
	hoverFlagsForTooltipMouse        ImGuiHoveredFlags
	hoverFlagsForTooltipNav          ImGuiHoveredFlags
}

struct ImGuiKeyData {
	down             bool
	downDuration     f32
	downDurationPrev f32
	analogValue      f32
}

struct ImVector_ImWchar {
	size     int
	capacity int
	data     &C.ImWchar
}

struct ImGuiIO {
	configFlags                                   ImGuiConfigFlags
	backendFlags                                  ImGuiBackendFlags
	displaySize                                   ImVec2
	deltaTime                                     f32
	iniSavingRate                                 f32
	iniFilename                                   &i8
	logFilename                                   &i8
	userData                                      voidptr
	fonts                                         &ImFontAtlas
	fontGlobalScale                               f32
	fontAllowUserScaling                          bool
	fontDefault                                   &ImFont
	displayFramebufferScale                       ImVec2
	configNavSwapGamepadButtons                   bool
	configNavMoveSetMousePos                      bool
	configNavCaptureKeyboard                      bool
	configNavEscapeClearFocusItem                 bool
	configNavEscapeClearFocusWindow               bool
	configNavCursorVisibleAuto                    bool
	configNavCursorVisibleAlways                  bool
	configDockingNoSplit                          bool
	configDockingWithShift                        bool
	configDockingAlwaysTabBar                     bool
	configDockingTransparentPayload               bool
	configViewportsNoAutoMerge                    bool
	configViewportsNoTaskBarIcon                  bool
	configViewportsNoDecoration                   bool
	configViewportsNoDefaultParent                bool
	mouseDrawCursor                               bool
	configMacOSXBehaviors                         bool
	configInputTrickleEventQueue                  bool
	configInputTextCursorBlink                    bool
	configInputTextEnterKeepActive                bool
	configDragClickToInputText                    bool
	configWindowsResizeFromEdges                  bool
	configWindowsMoveFromTitleBarOnly             bool
	configWindowsCopyContentsWithCtrlC            bool
	configScrollbarScrollByPage                   bool
	configMemoryCompactTimer                      f32
	mouseDoubleClickTime                          f32
	mouseDoubleClickMaxDist                       f32
	mouseDragThreshold                            f32
	keyRepeatDelay                                f32
	keyRepeatRate                                 f32
	configErrorRecovery                           bool
	configErrorRecoveryEnableAssert               bool
	configErrorRecoveryEnableDebugLog             bool
	configErrorRecoveryEnableTooltip              bool
	configDebugIsDebuggerPresent                  bool
	configDebugHighlightIdConflicts               bool
	configDebugHighlightIdConflictsShowItemPicker bool
	configDebugBeginReturnValueOnce               bool
	configDebugBeginReturnValueLoop               bool
	configDebugIgnoreFocusLoss                    bool
	configDebugIniSettings                        bool
	backendPlatformName                           &i8
	backendRendererName                           &i8
	backendPlatformUserData                       voidptr
	backendRendererUserData                       voidptr
	backendLanguageUserData                       voidptr
	wantCaptureMouse                              bool
	wantCaptureKeyboard                           bool
	wantTextInput                                 bool
	wantSetMousePos                               bool
	wantSaveIniSettings                           bool
	navActive                                     bool
	navVisible                                    bool
	framerate                                     f32
	metricsRenderVertices                         int
	metricsRenderIndices                          int
	metricsRenderWindows                          int
	metricsActiveWindows                          int
	mouseDelta                                    ImVec2
	ctx                                           &ImGuiContext
	mousePos                                      ImVec2
	mouseDown                                     [5]bool
	mouseWheel                                    f32
	mouseWheelH                                   f32
	mouseSource                                   ImGuiMouseSource
	mouseHoveredViewport                          ImGuiID
	keyCtrl                                       bool
	keyShift                                      bool
	keyAlt                                        bool
	keySuper                                      bool
	keyMods                                       ImGuiKeyChord
	keysData                                      [155]ImGuiKeyData
	wantCaptureMouseUnlessPopupClose              bool
	mousePosPrev                                  ImVec2
	mouseClickedPos                               [5]ImVec2
	mouseClickedTime                              [5]f64
	mouseClicked                                  [5]bool
	mouseDoubleClicked                            [5]bool
	mouseClickedCount                             [5]ImU16
	mouseClickedLastCount                         [5]ImU16
	mouseReleased                                 [5]bool
	mouseReleasedTime                             [5]f64
	mouseDownOwned                                [5]bool
	mouseDownOwnedUnlessPopupClose                [5]bool
	mouseWheelRequestAxisSwap                     bool
	mouseCtrlLeftAsRightClick                     bool
	mouseDownDuration                             [5]f32
	mouseDownDurationPrev                         [5]f32
	mouseDragMaxDistanceAbs                       [5]ImVec2
	mouseDragMaxDistanceSqr                       [5]f32
	penPressure                                   f32
	appFocusLost                                  bool
	appAcceptingEvents                            bool
	inputQueueSurrogate                           ImWchar16
	inputQueueCharacters                          ImVector_ImWchar
}

struct ImGuiInputTextCallbackData {
	ctx            &ImGuiContext
	eventFlag      ImGuiInputTextFlags
	flags          ImGuiInputTextFlags
	userData       voidptr
	eventChar      C.ImWchar
	eventKey       ImGuiKey
	buf            &i8
	bufTextLen     int
	bufSize        int
	bufDirty       bool
	cursorPos      int
	selectionStart int
	selectionEnd   int
}

struct ImGuiSizeCallbackData {
	userData    voidptr
	pos         ImVec2
	currentSize ImVec2
	desiredSize ImVec2
}

struct ImGuiWindowClass {
	classId                    ImGuiID
	parentViewportId           ImGuiID
	focusRouteParentWindowId   ImGuiID
	viewportFlagsOverrideSet   ImGuiViewportFlags
	viewportFlagsOverrideClear ImGuiViewportFlags
	tabItemFlagsOverrideSet    ImGuiTabItemFlags
	dockNodeFlagsOverrideSet   ImGuiDockNodeFlags
	dockingAlwaysTabBar        bool
	dockingAllowUnclassed      bool
}

struct ImGuiPayload {
	data           voidptr
	dataSize       int
	sourceId       ImGuiID
	sourceParentId ImGuiID
	dataFrameCount int
	dataType       [33]i8
	preview        bool
	delivery       bool
}

struct ImGuiOnceUponAFrame {
	refFrame int
}

struct ImGuiTextRange {
	b &i8
	e &i8
}

struct ImVector_ImGuiTextRange {
	size     int
	capacity int
	data     &ImGuiTextRange
}

struct ImVector_char {
	size     int
	capacity int
	data     &i8
}

struct ImGuiTextBuffer {
	buf ImVector_char
}

struct ImGuiStoragePair {
	key ImGuiID
}

struct ImVector_ImGuiStoragePair {
	size     int
	capacity int
	data     &ImGuiStoragePair
}

struct ImGuiStorage {
	data ImVector_ImGuiStoragePair
}

struct ImGuiListClipper {
	ctx              &ImGuiContext
	displayStart     int
	displayEnd       int
	itemsCount       int
	itemsHeight      f32
	startPosY        f32
	startSeekOffsetY f64
	tempData         voidptr
}

struct ImColor {
	value C.ImVec4
}

enum ImGuiMultiSelectFlags_ {
	none                      = 0
	single_select             = 1 << 0
	no_select_all             = 1 << 1
	no_range_select           = 1 << 2
	no_auto_select            = 1 << 3
	no_auto_clear             = 1 << 4
	no_auto_clear_on_reselect = 1 << 5
	box_select1d              = 1 << 6
	box_select2d              = 1 << 7
	box_select_no_scroll      = 1 << 8
	clear_on_escape           = 1 << 9
	clear_on_click_void       = 1 << 10
	scope_window              = 1 << 11
	scope_rect                = 1 << 12
	select_on_click           = 1 << 13
	select_on_click_release   = 1 << 14
	nav_wrap_x                = 1 << 16
}

struct ImVector_ImGuiSelectionRequest {
	size     int
	capacity int
	data     &ImGuiSelectionRequest
}

struct ImGuiMultiSelectIO {
	requests      ImVector_ImGuiSelectionRequest
	rangeSrcItem  ImGuiSelectionUserData
	navIdItem     ImGuiSelectionUserData
	navIdSelected bool
	rangeSrcReset bool
	itemsCount    int
}

enum ImGuiSelectionRequestType {
	none = 0
	set_all
	set_range
}

struct ImGuiSelectionRequest {
	type           ImGuiSelectionRequestType
	selected       bool
	rangeDirection ImS8
	rangeFirstItem ImGuiSelectionUserData
	rangeLastItem  ImGuiSelectionUserData
}

struct ImGuiSelectionBasicStorage {
	size                    int
	preserveOrder           bool
	userData                voidptr
	adapterIndexToStorageId fn (&ImGuiSelectionBasicStorage, int) ImGuiID
	_SelectionOrder         int
	_Storage                ImGuiStorage
}

struct ImDrawIdx {
	userData               voidptr
	adapterSetItemSelected fn (&C.ImGuiSelectionExternalStorage, int, bool)
}

type ImDrawCallback = fn (&ImDrawList, &ImDrawCmd)

struct ImDrawCmd {
	clipRect               C.ImVec4
	textureId              ImTextureID
	vtxOffset              u32
	idxOffset              u32
	elemCount              u32
	userCallback           ImDrawCallback
	userCallbackData       voidptr
	userCallbackDataSize   int
	userCallbackDataOffset int
}

struct ImDrawVert {
	pos ImVec2
	uv  ImVec2
	col ImU32
}

struct ImDrawCmdHeader {
	clipRect  C.ImVec4
	textureId ImTextureID
	vtxOffset u32
}

struct ImVector_ImDrawCmd {
	size     int
	capacity int
	data     &ImDrawCmd
}

struct ImVector_ImDrawIdx {
	size     int
	capacity int
	data     &ImDrawIdx
}

struct ImDrawChannel {
	_CmdBuffer ImVector_ImDrawCmd
	_IdxBuffer ImVector_ImDrawIdx
}

struct ImVector_ImDrawChannel {
	size     int
	capacity int
	data     &ImDrawChannel
}

struct ImDrawListSplitter {
	_Current  int
	_Count    int
	_Channels ImVector_ImDrawChannel
}

enum ImDrawFlags_ {
	none                       = 0
	closed                     = 1 << 0
	round_corners_top_left     = 1 << 4
	round_corners_top_right    = 1 << 5
	round_corners_bottom_left  = 1 << 6
	round_corners_bottom_right = 1 << 7
	round_corners_none         = 1 << 8
	round_corners_top          = 1 << 4 | 1 << 5
	round_corners_bottom       = 1 << 6 | 1 << 7
	round_corners_left         = 1 << 6 | 1 << 4
	round_corners_right        = 1 << 7 | 1 << 5
	round_corners_all          = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	round_corners_default_     = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	round_corners_mask_        = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8
}

enum ImDrawListFlags_ {
	none                       = 0
	anti_aliased_lines         = 1 << 0
	anti_aliased_lines_use_tex = 1 << 1
	anti_aliased_fill          = 1 << 2
	allow_vtx_offset           = 1 << 3
}

struct ImVector_ImDrawVert {
	size     int
	capacity int
	data     &ImDrawVert
}

struct ImVector_ImVec2 {
	size     int
	capacity int
	data     &ImVec2
}

struct ImVector_ImVec4 {
	size     int
	capacity int
	data     &C.ImVec4
}

struct ImVector_ImTextureID {
	size     int
	capacity int
	data     &ImTextureID
}

struct ImVector_ImU8 {
	size     int
	capacity int
	data     &ImU8
}

struct ImDrawList {
	cmdBuffer         ImVector_ImDrawCmd
	idxBuffer         ImVector_ImDrawIdx
	vtxBuffer         ImVector_ImDrawVert
	flags             ImDrawListFlags
	_VtxCurrentIdx    u32
	_Data             &ImDrawListSharedData
	_VtxWritePtr      &ImDrawVert
	_IdxWritePtr      &ImDrawIdx
	_Path             ImVector_ImVec2
	_CmdHeader        ImDrawCmdHeader
	_Splitter         ImDrawListSplitter
	_ClipRectStack    ImVector_ImVec4
	_TextureIdStack   ImVector_ImTextureID
	_CallbacksDataBuf ImVector_ImU8
	_FringeScale      f32
	_OwnerName        &i8
}

struct ImVector_ImDrawListPtr {
	size     int
	capacity int
	data     &&ImDrawList
}

struct ImDrawData {
	valid            bool
	cmdListsCount    int
	totalIdxCount    int
	totalVtxCount    int
	cmdLists         ImVector_ImDrawListPtr
	displayPos       ImVec2
	displaySize      ImVec2
	framebufferScale ImVec2
	ownerViewport    &ImGuiViewport
}

struct ImFontConfig {
	fontData             voidptr
	fontDataSize         int
	fontDataOwnedByAtlas bool
	mergeMode            bool
	pixelSnapH           bool
	fontNo               int
	oversampleH          int
	oversampleV          int
	sizePixels           f32
	glyphOffset          ImVec2
	glyphRanges          &C.ImWchar
	glyphMinAdvanceX     f32
	glyphMaxAdvanceX     f32
	glyphExtraAdvanceX   f32
	fontBuilderFlags     u32
	rasterizerMultiply   f32
	rasterizerDensity    f32
	ellipsisChar         C.ImWchar
	name                 [40]i8
	dstFont              &ImFont
}

struct ImFontGlyph {
	colored   u32
	visible   u32
	codepoint u32
	advanceX  f32
	x0        f32
	y0        f32
	x1        f32
	y1        f32
	u0        f32
	v0        f32
	u1        f32
	v1        f32
}

struct ImVector_ImU32 {
	size     int
	capacity int
	data     &ImU32
}

struct ImFontGlyphRangesBuilder {
	usedChars ImVector_ImU32
}

struct ImFontAtlasCustomRect {
	x             u16
	y             u16
	width         u16
	height        u16
	glyphID       u32
	glyphColored  u32
	glyphAdvanceX f32
	glyphOffset   ImVec2
	font          &ImFont
}

enum ImFontAtlasFlags_ {
	none                   = 0
	no_power_of_two_height = 1 << 0
	no_mouse_cursors       = 1 << 1
	no_baked_lines         = 1 << 2
}

struct ImVector_ImFontPtr {
	size     int
	capacity int
	data     &&ImFont
}

struct ImVector_ImFontAtlasCustomRect {
	size     int
	capacity int
	data     &ImFontAtlasCustomRect
}

struct ImVector_ImFontConfig {
	size     int
	capacity int
	data     &ImFontConfig
}

struct ImFontAtlas {
	flags              ImFontAtlasFlags
	texID              ImTextureID
	texDesiredWidth    int
	texGlyphPadding    int
	userData           voidptr
	locked             bool
	texReady           bool
	texPixelsUseColors bool
	texPixelsAlpha8    &u8
	texPixelsRGBA32    &u32
	texWidth           int
	texHeight          int
	texUvScale         ImVec2
	texUvWhitePixel    ImVec2
	fonts              ImVector_ImFontPtr
	customRects        ImVector_ImFontAtlasCustomRect
	sources            ImVector_ImFontConfig
	texUvLines         [33]C.ImVec4
	fontBuilderIO      &ImFontBuilderIO
	fontBuilderFlags   u32
	packIdMouseCursors int
	packIdLines        int
}

struct ImVector_float {
	size     int
	capacity int
	data     &f32
}

struct ImVector_ImU16 {
	size     int
	capacity int
	data     &ImU16
}

struct ImVector_ImFontGlyph {
	size     int
	capacity int
	data     &ImFontGlyph
}

struct ImFont {
	indexAdvanceX       ImVector_float
	fallbackAdvanceX    f32
	fontSize            f32
	indexLookup         ImVector_ImU16
	glyphs              ImVector_ImFontGlyph
	fallbackGlyph       &ImFontGlyph
	containerAtlas      &ImFontAtlas
	sources             &ImFontConfig
	sourcesCount        i16
	ellipsisCharCount   i16
	ellipsisChar        C.ImWchar
	fallbackChar        C.ImWchar
	ellipsisWidth       f32
	ellipsisCharStep    f32
	scale               f32
	ascent              f32
	descent             f32
	metricsTotalSurface int
	dirtyLookupTables   bool
	used8kPagesMap      [17]ImU8
}

enum ImGuiViewportFlags_ {
	none                   = 0
	is_platform_window     = 1 << 0
	is_platform_monitor    = 1 << 1
	owned_by_app           = 1 << 2
	no_decoration          = 1 << 3
	no_task_bar_icon       = 1 << 4
	no_focus_on_appearing  = 1 << 5
	no_focus_on_click      = 1 << 6
	no_inputs              = 1 << 7
	no_renderer_clear      = 1 << 8
	no_auto_merge          = 1 << 9
	top_most               = 1 << 10
	can_host_other_windows = 1 << 11
	is_minimized           = 1 << 12
	is_focused             = 1 << 13
}

struct ImGuiViewport {
	iD                    ImGuiID
	flags                 ImGuiViewportFlags
	pos                   ImVec2
	size                  ImVec2
	workPos               ImVec2
	workSize              ImVec2
	dpiScale              f32
	parentViewportId      ImGuiID
	drawData              &ImDrawData
	rendererUserData      voidptr
	platformUserData      voidptr
	platformHandle        voidptr
	platformHandleRaw     voidptr
	platformWindowCreated bool
	platformRequestMove   bool
	platformRequestResize bool
	platformRequestClose  bool
}

struct ImVector_ImGuiPlatformMonitor {
	size     int
	capacity int
	data     &ImGuiPlatformMonitor
}

struct ImVector_ImGuiViewportPtr {
	size     int
	capacity int
	data     &&ImGuiViewport
}

struct ImGuiPlatformIO {
	platform_GetClipboardTextFn      fn (&ImGuiContext) &i8
	platform_SetClipboardTextFn      fn (&ImGuiContext, &i8)
	platform_ClipboardUserData       voidptr
	platform_OpenInShellFn           fn (&ImGuiContext, &i8) bool
	platform_OpenInShellUserData     voidptr
	platform_SetImeDataFn            fn (&ImGuiContext, &ImGuiViewport, &ImGuiPlatformImeData)
	platform_ImeUserData             voidptr
	platform_LocaleDecimalPoint      C.ImWchar
	renderer_RenderState             voidptr
	platform_CreateWindow            fn (&ImGuiViewport)
	platform_DestroyWindow           fn (&ImGuiViewport)
	platform_ShowWindow              fn (&ImGuiViewport)
	platform_SetWindowPos            fn (&ImGuiViewport, ImVec2)
	platform_GetWindowPos            fn (&ImGuiViewport) ImVec2
	platform_SetWindowSize           fn (&ImGuiViewport, ImVec2)
	platform_GetWindowSize           fn (&ImGuiViewport) ImVec2
	platform_SetWindowFocus          fn (&ImGuiViewport)
	platform_GetWindowFocus          fn (&ImGuiViewport) bool
	platform_GetWindowMinimized      fn (&ImGuiViewport) bool
	platform_SetWindowTitle          fn (&ImGuiViewport, &i8)
	platform_SetWindowAlpha          fn (&ImGuiViewport, f32)
	platform_UpdateWindow            fn (&ImGuiViewport)
	platform_RenderWindow            fn (&ImGuiViewport, voidptr)
	platform_SwapBuffers             fn (&ImGuiViewport, voidptr)
	platform_GetWindowDpiScale       fn (&ImGuiViewport) f32
	platform_OnChangedViewport       fn (&ImGuiViewport)
	platform_GetWindowWorkAreaInsets fn (&ImGuiViewport) C.ImVec4
	platform_CreateVkSurface         fn (&ImGuiViewport, ImU64, voidptr, &ImU64) int
	renderer_CreateWindow            fn (&ImGuiViewport)
	renderer_DestroyWindow           fn (&ImGuiViewport)
	renderer_SetWindowSize           fn (&ImGuiViewport, ImVec2)
	renderer_RenderWindow            fn (&ImGuiViewport, voidptr)
	renderer_SwapBuffers             fn (&ImGuiViewport, voidptr)
	monitors                         ImVector_ImGuiPlatformMonitor
	viewports                        ImVector_ImGuiViewportPtr
}

struct ImGuiPlatformMonitor {
	mainPos        ImVec2
	mainSize       ImVec2
	workPos        ImVec2
	workSize       ImVec2
	dpiScale       f32
	platformHandle voidptr
}

struct ImGuiPlatformImeData {
	wantVisible     bool
	inputPos        ImVec2
	inputLineHeight f32
}

type ImGuiDataAuthority = int
type ImGuiLayoutType = int
type ImGuiActivateFlags = int
type ImGuiDebugLogFlags = int
type ImGuiFocusRequestFlags = int
type ImGuiItemStatusFlags = int
type ImGuiOldColumnFlags = int
type ImGuiLogFlags = int
type ImGuiNavRenderCursorFlags = int
type ImGuiNavMoveFlags = int
type ImGuiNextItemDataFlags = int
type ImGuiNextWindowDataFlags = int
type ImGuiScrollFlags = int
type ImGuiSeparatorFlags = int
type ImGuiTextFlags = int
type ImGuiTooltipFlags = int
type ImGuiTypingSelectFlags = int
type ImGuiWindowRefreshFlags = int
type ImFileHandle = &C.FILE

struct ImVec1 {
	x f32
}

struct ImVec2ih {
	x i16
	y i16
}

struct ImBitArrayPtr {
	min ImVec2
	max ImVec2
}

struct ImPoolIdx {
	storage ImVector_ImU32
}

struct ImVector_int {
	size     int
	capacity int
	data     &int
}

struct ImGuiTextIndex {
	lineOffsets ImVector_int
	endOffset   int
}

struct ImDrawListSharedData {
	texUvWhitePixel       ImVec2
	texUvLines            &C.ImVec4
	font                  &ImFont
	fontSize              f32
	fontScale             f32
	curveTessellationTol  f32
	circleSegmentMaxError f32
	initialFringeScale    f32
	initialFlags          ImDrawListFlags
	clipRectFullscreen    C.ImVec4
	tempBuffer            ImVector_ImVec2
	arcFastVtx            [48]ImVec2
	arcFastRadiusCutoff   f32
	circleSegmentCounts   [64]ImU8
}

struct ImDrawDataBuilder {
	layers     [2]&ImVector_ImDrawListPtr
	layerData1 ImVector_ImDrawListPtr
}

struct ImGuiStyleVarInfo {
	count    ImU32
	dataType ImGuiDataType
	offset   ImU32
}

struct ImGuiColorMod {
	col         ImGuiCol
	backupValue C.ImVec4
}

struct ImGuiStyleMod {
	varIdx ImGuiStyleVar
}

struct ImGuiDataTypeStorage {
	data [8]ImU8
}

struct ImGuiDataTypeInfo {
	size     usize
	name     &i8
	printFmt &i8
	scanFmt  &i8
}

enum ImGuiDataTypePrivate_ {
	pointer = int(ImGuiDataType_.count)
	id
}

enum ImGuiItemFlagsPrivate_ {
	disabled                   = 1 << 10
	read_only                  = 1 << 11
	mixed_value                = 1 << 12
	no_window_hoverable_check  = 1 << 13
	allow_overlap              = 1 << 14
	no_nav_disable_mouse_hover = 1 << 15
	no_mark_edited             = 1 << 16
	inputable                  = 1 << 20
	has_selection_user_data    = 1 << 21
	is_multi_select            = 1 << 22
	default_                   = 1 << 4
}

enum ImGuiItemStatusFlags_ {
	none              = 0
	hovered_rect      = 1 << 0
	has_display_rect  = 1 << 1
	edited            = 1 << 2
	toggled_selection = 1 << 3
	toggled_open      = 1 << 4
	has_deactivated   = 1 << 5
	deactivated       = 1 << 6
	hovered_window    = 1 << 7
	visible           = 1 << 8
	has_clip_rect     = 1 << 9
	has_shortcut      = 1 << 10
}

enum ImGuiHoveredFlagsPrivate_ {
	delay_mask_                        = 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
	allowed_mask_for_is_window_hovered = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 7 | 1 << 12 | 1 << 13
	allowed_mask_for_is_item_hovered   = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
}

enum ImGuiInputTextFlagsPrivate_ {
	multiline              = 1 << 26
	merged_item            = 1 << 27
	localize_decimal_point = 1 << 28
}

enum ImGuiButtonFlagsPrivate_ {
	pressed_on_click                  = 1 << 4
	pressed_on_click_release          = 1 << 5
	pressed_on_click_release_anywhere = 1 << 6
	pressed_on_release                = 1 << 7
	pressed_on_double_click           = 1 << 8
	pressed_on_drag_drop_hold         = 1 << 9
	flatten_children                  = 1 << 11
	allow_overlap                     = 1 << 12
	align_text_base_line              = 1 << 15
	no_key_mods_allowed               = 1 << 16
	no_holding_active_id              = 1 << 17
	no_nav_focus                      = 1 << 18
	no_hovered_on_focus               = 1 << 19
	no_set_key_owner                  = 1 << 20
	no_test_key_owner                 = 1 << 21
	pressed_on_mask_                  = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8 | 1 << 9
	pressed_on_default_               = 1 << 5
}

enum ImGuiComboFlagsPrivate_ {
	custom_preview = 1 << 20
}

enum ImGuiSliderFlagsPrivate_ {
	vertical  = 1 << 20
	read_only = 1 << 21
}

enum ImGuiSelectableFlagsPrivate_ {
	no_holding_active_id     = 1 << 20
	select_on_nav            = 1 << 21
	select_on_click          = 1 << 22
	select_on_release        = 1 << 23
	span_avail_width         = 1 << 24
	set_nav_id_on_hover      = 1 << 25
	no_pad_with_half_spacing = 1 << 26
	no_set_key_owner         = 1 << 27
}

enum ImGuiTreeNodeFlagsPrivate_ {
	clip_label_for_trailing_button = 1 << 28
	upside_down_arrow              = 1 << 29
	open_on_mask_                  = 1 << 6 | 1 << 7
}

enum ImGuiSeparatorFlags_ {
	none             = 0
	horizontal       = 1 << 0
	vertical         = 1 << 1
	span_all_columns = 1 << 2
}

enum ImGuiFocusRequestFlags_ {
	none                  = 0
	restore_focused_child = 1 << 0
	unless_below_modal    = 1 << 1
}

enum ImGuiTextFlags_ {
	none                            = 0
	no_width_for_large_clipped_text = 1 << 0
}

enum ImGuiTooltipFlags_ {
	none              = 0
	override_previous = 1 << 1
}

enum ImGuiLayoutType_ {
	horizontal = 0
	vertical   = 1
}

enum ImGuiLogFlags_ {
	none             = 0
	output_tty       = 1 << 0
	output_file      = 1 << 1
	output_buffer    = 1 << 2
	output_clipboard = 1 << 3
	output_mask_     = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
}

enum ImGuiAxis {
	none = -1
	x    = 0
	y    = 1
}

enum ImGuiPlotType {
	lines
	histogram
}

struct ImGuiComboPreviewData {
	previewRect                  C.ImRect
	backupCursorPos              ImVec2
	backupCursorMaxPos           ImVec2
	backupCursorPosPrevLine      ImVec2
	backupPrevLineTextBaseOffset f32
	backupLayout                 ImGuiLayoutType
}

struct ImGuiGroupData {
	windowID                     ImGuiID
	backupCursorPos              ImVec2
	backupCursorMaxPos           ImVec2
	backupCursorPosPrevLine      ImVec2
	backupIndent                 ImVec1
	backupGroupOffset            ImVec1
	backupCurrLineSize           ImVec2
	backupCurrLineTextBaseOffset f32
	backupActiveIdIsAlive        ImGuiID
	backupDeactivatedIdIsAlive   bool
	backupHoveredIdIsAlive       bool
	backupIsSameLine             bool
	emitItem                     bool
}

struct ImGuiMenuColumns {
	totalWidth     ImU32
	nextTotalWidth ImU32
	spacing        ImU16
	offsetIcon     ImU16
	offsetLabel    ImU16
	offsetShortcut ImU16
	offsetMark     ImU16
	widths         [4]ImU16
}

struct ImGuiInputTextDeactivatedState {
	iD    ImGuiID
	textA ImVector_char
}

type ImStbTexteditState = voidptr

struct ImGuiInputTextState {
	ctx                  &ImGuiContext
	stb                  &ImStbTexteditState
	flags                ImGuiInputTextFlags
	iD                   ImGuiID
	textLen              int
	textSrc              &i8
	textA                ImVector_char
	textToRevertTo       ImVector_char
	callbackTextBackup   ImVector_char
	bufCapacity          int
	scroll               ImVec2
	cursorAnim           f32
	cursorFollow         bool
	selectedAllMouseLock bool
	edited               bool
	wantReloadUserBuf    bool
	reloadSelectionStart int
	reloadSelectionEnd   int
}

enum ImGuiWindowRefreshFlags_ {
	none                 = 0
	try_to_avoid_refresh = 1 << 0
	refresh_on_hover     = 1 << 1
	refresh_on_focus     = 1 << 2
}

enum ImGuiNextWindowDataFlags_ {
	none                = 0
	has_pos             = 1 << 0
	has_size            = 1 << 1
	has_content_size    = 1 << 2
	has_collapsed       = 1 << 3
	has_size_constraint = 1 << 4
	has_focus           = 1 << 5
	has_bg_alpha        = 1 << 6
	has_scroll          = 1 << 7
	has_window_flags    = 1 << 8
	has_child_flags     = 1 << 9
	has_refresh_policy  = 1 << 10
	has_viewport        = 1 << 11
	has_dock            = 1 << 12
	has_window_class    = 1 << 13
}

struct ImGuiNextWindowData {
	hasFlags             ImGuiNextWindowDataFlags
	posCond              ImGuiCond
	sizeCond             ImGuiCond
	collapsedCond        ImGuiCond
	dockCond             ImGuiCond
	posVal               ImVec2
	posPivotVal          ImVec2
	sizeVal              ImVec2
	contentSizeVal       ImVec2
	scrollVal            ImVec2
	windowFlags          ImGuiWindowFlags
	childFlags           ImGuiChildFlags
	posUndock            bool
	collapsedVal         bool
	sizeConstraintRect   C.ImRect
	sizeCallback         C.ImGuiSizeCallback
	sizeCallbackUserData voidptr
	bgAlphaVal           f32
	viewportId           ImGuiID
	dockId               ImGuiID
	windowClass          ImGuiWindowClass
	menuBarOffsetMinVal  ImVec2
	refreshFlagsVal      ImGuiWindowRefreshFlags
}

enum ImGuiNextItemDataFlags_ {
	none           = 0
	has_width      = 1 << 0
	has_open       = 1 << 1
	has_shortcut   = 1 << 2
	has_ref_val    = 1 << 3
	has_storage_id = 1 << 4
}

struct ImGuiNextItemData {
	hasFlags          ImGuiNextItemDataFlags
	itemFlags         ImGuiItemFlags
	focusScopeId      ImGuiID
	selectionUserData ImGuiSelectionUserData
	width             f32
	shortcut          ImGuiKeyChord
	shortcutFlags     ImGuiInputFlags
	openVal           bool
	openCond          ImU8
	refVal            ImGuiDataTypeStorage
	storageId         ImGuiID
}

struct ImGuiLastItemData {
	iD          ImGuiID
	itemFlags   ImGuiItemFlags
	statusFlags ImGuiItemStatusFlags
	rect        C.ImRect
	navRect     C.ImRect
	displayRect C.ImRect
	clipRect    C.ImRect
	shortcut    ImGuiKeyChord
}

struct ImGuiTreeNodeStackData {
	iD        ImGuiID
	treeFlags ImGuiTreeNodeFlags
	itemFlags ImGuiItemFlags
	navRect   C.ImRect
}

struct ImGuiErrorRecoveryState {
	sizeOfWindowStack     i16
	sizeOfIDStack         i16
	sizeOfTreeStack       i16
	sizeOfColorStack      i16
	sizeOfStyleVarStack   i16
	sizeOfFontStack       i16
	sizeOfFocusScopeStack i16
	sizeOfGroupStack      i16
	sizeOfItemFlagsStack  i16
	sizeOfBeginPopupStack i16
	sizeOfDisabledStack   i16
}

struct ImGuiWindowStackData {
	window                              &ImGuiWindow
	parentLastItemDataBackup            ImGuiLastItemData
	stackSizesInBegin                   ImGuiErrorRecoveryState
	disabledOverrideReenable            bool
	disabledOverrideReenableAlphaBackup f32
}

struct ImGuiShrinkWidthItem {
	index        int
	width        f32
	initialWidth f32
}

struct ImGuiPtrOrIndex {
	ptr   voidptr
	index int
}

struct ImGuiDeactivatedItemData {
	iD                  ImGuiID
	elapseFrame         int
	hasBeenEditedBefore bool
	isAlive             bool
}

enum ImGuiPopupPositionPolicy {
	default
	combo_box
	tooltip
}

struct ImGuiPopupData {
	popupId          ImGuiID
	window           &ImGuiWindow
	restoreNavWindow &ImGuiWindow
	parentNavLayer   int
	openFrameCount   int
	openParentId     ImGuiID
	openPopupPos     ImVec2
	openMousePos     ImVec2
}

struct ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN {
	storage [5]ImU32
}

type ImBitArrayForNamedKeys = ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN

enum ImGuiInputEventType {
	none = 0
	mouse_pos
	mouse_wheel
	mouse_button
	mouse_viewport
	key
	text
	focus
	count
}

enum ImGuiInputSource {
	none = 0
	mouse
	keyboard
	gamepad
	count
}

struct ImGuiInputEventMousePos {
	posX        f32
	posY        f32
	mouseSource ImGuiMouseSource
}

struct ImGuiInputEventMouseWheel {
	wheelX      f32
	wheelY      f32
	mouseSource ImGuiMouseSource
}

struct ImGuiInputEventMouseButton {
	button      int
	down        bool
	mouseSource ImGuiMouseSource
}

struct ImGuiInputEventMouseViewport {
	hoveredViewportID ImGuiID
}

struct ImGuiInputEventKey {
	key         ImGuiKey
	down        bool
	analogValue f32
}

struct ImGuiInputEventText {
	char u32
}

struct ImGuiInputEventAppFocused {
	focused bool
}

struct ImGuiKeyRoutingIndex {
	type              ImGuiInputEventType
	source            ImGuiInputSource
	eventId           ImU32
	addedByTestEngine bool
}

struct ImGuiKeyRoutingData {
	nextEntryIndex   ImGuiKeyRoutingIndex
	mods             ImU16
	routingCurrScore ImU8
	routingNextScore ImU8
	routingCurr      ImGuiID
	routingNext      ImGuiID
}

struct ImVector_ImGuiKeyRoutingData {
	size     int
	capacity int
	data     &ImGuiKeyRoutingData
}

struct ImGuiKeyRoutingTable {
	index       [155]ImGuiKeyRoutingIndex
	entries     ImVector_ImGuiKeyRoutingData
	entriesNext ImVector_ImGuiKeyRoutingData
}

struct ImGuiKeyOwnerData {
	ownerCurr        ImGuiID
	ownerNext        ImGuiID
	lockThisFrame    bool
	lockUntilRelease bool
}

enum ImGuiInputFlagsPrivate_ {
	repeat_rate_default                    = 1 << 1
	repeat_rate_nav_move                   = 1 << 2
	repeat_rate_nav_tweak                  = 1 << 3
	repeat_until_release                   = 1 << 4
	repeat_until_key_mods_change           = 1 << 5
	repeat_until_key_mods_change_from_none = 1 << 6
	repeat_until_other_key_press           = 1 << 7
	lock_this_frame                        = 1 << 20
	lock_until_release                     = 1 << 21
	cond_hovered                           = 1 << 22
	cond_active                            = 1 << 23
	cond_default_                          = 1 << 22 | 1 << 23
	repeat_rate_mask_                      = 1 << 1 | 1 << 2 | 1 << 3
	repeat_until_mask_                     = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	repeat_mask_                           = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	cond_mask_                             = 1 << 22 | 1 << 23
	route_type_mask_                       = 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13
	route_options_mask_                    = 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
	supported_by_is_key_pressed            = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	supported_by_is_mouse_clicked          = 1 << 0
	supported_by_shortcut                  = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
	supported_by_set_next_item_shortcut    = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17 | 1 << 18
	supported_by_set_key_owner             = 1 << 20 | 1 << 21
	supported_by_set_item_key_owner        = 1 << 20 | 1 << 21 | 1 << 22 | 1 << 23
}

struct ImGuiListClipperRange {
	min                 int
	max                 int
	posToIndexConvert   bool
	posToIndexOffsetMin ImS8
	posToIndexOffsetMax ImS8
}

struct ImVector_ImGuiListClipperRange {
	size     int
	capacity int
	data     &ImGuiListClipperRange
}

struct ImGuiListClipperData {
	listClipper     &ImGuiListClipper
	lossynessOffset f32
	stepNo          int
	itemsFrozen     int
	ranges          ImVector_ImGuiListClipperRange
}

enum ImGuiActivateFlags_ {
	none                  = 0
	prefer_input          = 1 << 0
	prefer_tweak          = 1 << 1
	try_to_preserve_state = 1 << 2
	from_tabbing          = 1 << 3
	from_shortcut         = 1 << 4
}

enum ImGuiScrollFlags_ {
	none                  = 0
	keep_visible_edge_x   = 1 << 0
	keep_visible_edge_y   = 1 << 1
	keep_visible_center_x = 1 << 2
	keep_visible_center_y = 1 << 3
	always_center_x       = 1 << 4
	always_center_y       = 1 << 5
	no_scroll_parent      = 1 << 6
	mask_x_               = 1 << 0 | 1 << 2 | 1 << 4
	mask_y_               = 1 << 1 | 1 << 3 | 1 << 5
}

enum ImGuiNavRenderCursorFlags_ {
	none        = 0
	compact     = 1 << 1
	always_draw = 1 << 2
	no_rounding = 1 << 3
}

enum ImGuiNavMoveFlags_ {
	none                      = 0
	loop_x                    = 1 << 0
	loop_y                    = 1 << 1
	wrap_x                    = 1 << 2
	wrap_y                    = 1 << 3
	wrap_mask_                = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
	allow_current_nav_id      = 1 << 4
	also_score_visible_set    = 1 << 5
	scroll_to_edge_y          = 1 << 6
	forwarded                 = 1 << 7
	debug_no_result           = 1 << 8
	focus_api                 = 1 << 9
	is_tabbing                = 1 << 10
	is_page_move              = 1 << 11
	activate                  = 1 << 12
	no_select                 = 1 << 13
	no_set_nav_cursor_visible = 1 << 14
	no_clear_active_id        = 1 << 15
}

enum ImGuiNavLayer {
	main = 0
	menu = 1
	count
}

struct ImGuiNavItemData {
	window            &ImGuiWindow
	iD                ImGuiID
	focusScopeId      ImGuiID
	rectRel           C.ImRect
	itemFlags         ImGuiItemFlags
	distBox           f32
	distCenter        f32
	distAxial         f32
	selectionUserData ImGuiSelectionUserData
}

struct ImGuiFocusScopeData {
	iD       ImGuiID
	windowID ImGuiID
}

enum ImGuiTypingSelectFlags_ {
	none                   = 0
	allow_backspace        = 1 << 0
	allow_single_char_mode = 1 << 1
}

struct ImGuiTypingSelectRequest {
	flags           ImGuiTypingSelectFlags
	searchBufferLen int
	searchBuffer    &i8
	selectRequest   bool
	singleCharMode  bool
	singleCharSize  ImS8
}

struct ImGuiTypingSelectState {
	request            ImGuiTypingSelectRequest
	searchBuffer       [64]i8
	focusScope         ImGuiID
	lastRequestFrame   int
	lastRequestTime    f32
	singleCharModeLock bool
}

enum ImGuiOldColumnFlags_ {
	none                      = 0
	no_border                 = 1 << 0
	no_resize                 = 1 << 1
	no_preserve_widths        = 1 << 2
	no_force_within_window    = 1 << 3
	grow_parent_contents_size = 1 << 4
}

struct ImGuiOldColumnData {
	offsetNorm             f32
	offsetNormBeforeResize f32
	flags                  ImGuiOldColumnFlags
	clipRect               C.ImRect
}

struct ImVector_ImGuiOldColumnData {
	size     int
	capacity int
	data     &ImGuiOldColumnData
}

struct ImGuiOldColumns {
	iD                       ImGuiID
	flags                    ImGuiOldColumnFlags
	isFirstFrame             bool
	isBeingResized           bool
	current                  int
	count                    int
	offMinX                  f32
	offMaxX                  f32
	lineMinY                 f32
	lineMaxY                 f32
	hostCursorPosY           f32
	hostCursorMaxPosX        f32
	hostInitialClipRect      C.ImRect
	hostBackupClipRect       C.ImRect
	hostBackupParentWorkRect C.ImRect
	columns                  ImVector_ImGuiOldColumnData
	splitter                 ImDrawListSplitter
}

struct ImGuiBoxSelectState {
	iD                    ImGuiID
	isActive              bool
	isStarting            bool
	isStartedFromVoid     bool
	isStartedSetNavIdOnce bool
	requestClear          bool
	keyMods               ImGuiKeyChord
	startPosRel           ImVec2
	endPosRel             ImVec2
	scrollAccum           ImVec2
	window                &ImGuiWindow
	unclipMode            bool
	unclipRect            C.ImRect
	boxSelectRectPrev     C.ImRect
	boxSelectRectCurr     C.ImRect
}

struct ImGuiMultiSelectTempData {
	iO                 ImGuiMultiSelectIO
	storage            &ImGuiMultiSelectState
	focusScopeId       ImGuiID
	flags              ImGuiMultiSelectFlags
	scopeRectMin       ImVec2
	backupCursorMaxPos ImVec2
	lastSubmittedItem  ImGuiSelectionUserData
	boxSelectId        ImGuiID
	keyMods            ImGuiKeyChord
	loopRequestSetAll  ImS8
	isEndIO            bool
	isFocused          bool
	isKeyboardSetRange bool
	navIdPassedBy      bool
	rangeSrcPassedBy   bool
	rangeDstPassedBy   bool
}

struct ImGuiMultiSelectState {
	window            &ImGuiWindow
	iD                ImGuiID
	lastFrameActive   int
	lastSelectionSize int
	rangeSelected     ImS8
	navIdSelected     ImS8
	rangeSrcItem      ImGuiSelectionUserData
	navIdItem         ImGuiSelectionUserData
}

enum ImGuiDockNodeFlagsPrivate_ {
	dock_space                    = 1 << 10
	central_node                  = 1 << 11
	no_tab_bar                    = 1 << 12
	hidden_tab_bar                = 1 << 13
	no_window_menu_button         = 1 << 14
	no_close_button               = 1 << 15
	no_resize_x                   = 1 << 16
	no_resize_y                   = 1 << 17
	docked_windows_in_focus_route = 1 << 18
	no_docking_split_other        = 1 << 19
	no_docking_over_me            = 1 << 20
	no_docking_over_other         = 1 << 21
	no_docking_over_empty         = 1 << 22
	no_docking                    = 1 << 20 | 1 << 21 | 1 << 22 | 1 << 4 | 1 << 19
	shared_flags_inherit_mask_    = int(~0)
	no_resize_flags_mask_         = 1 << 5 | 1 << 16 | 1 << 17
	local_flags_transfer_mask_    = 1 << 4 | 1 << 5 | 1 << 16 | 1 << 17 | 1 << 6 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15
	saved_flags_mask_             = 1 << 5 | 1 << 16 | 1 << 17 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15
}

enum ImGuiDataAuthority_ {
	auto
	dock_node
	window
}

enum ImGuiDockNodeState {
	unknown
	host_window_hidden_because_single_window
	host_window_hidden_because_windows_are_resizing
	host_window_visible
}

struct ImVector_ImGuiWindowPtr {
	size     int
	capacity int
	data     &&ImGuiWindow
}

struct ImGuiDockNode {
	iD                     ImGuiID
	sharedFlags            ImGuiDockNodeFlags
	localFlags             ImGuiDockNodeFlags
	localFlagsInWindows    ImGuiDockNodeFlags
	mergedFlags            ImGuiDockNodeFlags
	state                  ImGuiDockNodeState
	parentNode             &ImGuiDockNode
	childNodes             [2]&ImGuiDockNode
	windows                ImVector_ImGuiWindowPtr
	tabBar                 &C.ImGuiTabBar
	pos                    ImVec2
	size                   ImVec2
	sizeRef                ImVec2
	splitAxis              ImGuiAxis
	windowClass            ImGuiWindowClass
	lastBgColor            ImU32
	hostWindow             &ImGuiWindow
	visibleWindow          &ImGuiWindow
	centralNode            &ImGuiDockNode
	onlyNodeWithWindows    &ImGuiDockNode
	countNodeWithWindows   int
	lastFrameAlive         int
	lastFrameActive        int
	lastFrameFocused       int
	lastFocusedNodeId      ImGuiID
	selectedTabId          ImGuiID
	wantCloseTabId         ImGuiID
	refViewportId          ImGuiID
	authorityForPos        ImGuiDataAuthority
	authorityForSize       ImGuiDataAuthority
	authorityForViewport   ImGuiDataAuthority
	isVisible              bool
	isFocused              bool
	isBgDrawnThisFrame     bool
	hasCloseButton         bool
	hasWindowMenuButton    bool
	hasCentralNodeChild    bool
	wantCloseAll           bool
	wantLockSizeOnce       bool
	wantMouseMove          bool
	wantHiddenTabBarUpdate bool
	wantHiddenTabBarToggle bool
}

enum ImGuiWindowDockStyleCol {
	text
	tab_hovered
	tab_focused
	tab_selected
	tab_selected_overline
	tab_dimmed
	tab_dimmed_selected
	tab_dimmed_selected_overline
	count
}

struct ImGuiWindowDockStyle {
	colors [8]ImU32
}

struct ImVector_ImGuiDockRequest {
	size     int
	capacity int
	data     &C.ImGuiDockRequest
}

struct ImVector_ImGuiDockNodeSettings {
	size     int
	capacity int
	data     &C.ImGuiDockNodeSettings
}

struct ImGuiDockContext {
	nodes           ImGuiStorage
	requests        ImVector_ImGuiDockRequest
	nodesSettings   ImVector_ImGuiDockNodeSettings
	wantFullRebuild bool
}

struct ImGuiViewportP {
	_ImGuiViewport          ImGuiViewport
	window                  &ImGuiWindow
	idx                     int
	lastFrameActive         int
	lastFocusedStampCount   int
	lastNameHash            ImGuiID
	lastPos                 ImVec2
	lastSize                ImVec2
	alpha                   f32
	lastAlpha               f32
	lastFocusedHadNavWindow bool
	platformMonitor         i16
	bgFgDrawListsLastFrame  [2]int
	bgFgDrawLists           [2]&ImDrawList
	drawDataP               ImDrawData
	drawDataBuilder         ImDrawDataBuilder
	lastPlatformPos         ImVec2
	lastPlatformSize        ImVec2
	lastRendererSize        ImVec2
	workInsetMin            ImVec2
	workInsetMax            ImVec2
	buildWorkInsetMin       ImVec2
	buildWorkInsetMax       ImVec2
}

struct ImGuiWindowSettings {
	iD          ImGuiID
	pos         ImVec2ih
	size        ImVec2ih
	viewportPos ImVec2ih
	viewportId  ImGuiID
	dockId      ImGuiID
	classId     ImGuiID
	dockOrder   i16
	collapsed   bool
	isChild     bool
	wantApply   bool
	wantDelete  bool
}

struct ImGuiSettingsHandler {
	typeName   &i8
	typeHash   ImGuiID
	clearAllFn fn (&ImGuiContext, &ImGuiSettingsHandler)
	readInitFn fn (&ImGuiContext, &ImGuiSettingsHandler)
	readOpenFn fn (&ImGuiContext, &ImGuiSettingsHandler, &i8) voidptr
	readLineFn fn (&ImGuiContext, &ImGuiSettingsHandler, voidptr, &i8)
	applyAllFn fn (&ImGuiContext, &ImGuiSettingsHandler)
	writeAllFn fn (&ImGuiContext, &ImGuiSettingsHandler, &ImGuiTextBuffer)
	userData   voidptr
}

enum ImGuiLocKey {
	version_str                         = 0
	table_size_one                      = 1
	table_size_all_fit                  = 2
	table_size_all_default              = 3
	table_reset_order                   = 4
	windowing_main_menu_bar             = 5
	windowing_popup                     = 6
	windowing_untitled                  = 7
	open_link_s                         = 8
	copy_link                           = 9
	docking_hide_tab_bar                = 10
	docking_hold_shift_to_dock          = 11
	docking_drag_to_undock_or_move_node = 12
	count                               = 13
}

struct ImGuiErrorCallback {
	key  ImGuiLocKey
	text &i8
}

enum ImGuiDebugLogFlags_ {
	none                  = 0
	event_error           = 1 << 0
	event_active_id       = 1 << 1
	event_focus           = 1 << 2
	event_popup           = 1 << 3
	event_nav             = 1 << 4
	event_clipper         = 1 << 5
	event_selection       = 1 << 6
	event_io              = 1 << 7
	event_font            = 1 << 8
	event_input_routing   = 1 << 9
	event_docking         = 1 << 10
	event_viewport        = 1 << 11
	event_mask_           = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8 | 1 << 9 | 1 << 10 | 1 << 11
	output_to_tty         = 1 << 20
	output_to_test_engine = 1 << 21
}

struct ImGuiDebugAllocEntry {
	frameCount int
	allocCount ImS16
	freeCount  ImS16
}

struct ImGuiDebugAllocInfo {
	totalAllocCount int
	totalFreeCount  int
	lastEntriesIdx  ImS16
	lastEntriesBuf  [6]ImGuiDebugAllocEntry
}

struct ImGuiMetricsConfig {
	showDebugLog             bool
	showIDStackTool          bool
	showWindowsRects         bool
	showWindowsBeginOrder    bool
	showTablesRects          bool
	showDrawCmdMesh          bool
	showDrawCmdBoundingBoxes bool
	showTextEncodingViewer   bool
	showDockingNodes         bool
	showWindowsRectsType     int
	showTablesRectsType      int
	highlightMonitorIdx      int
	highlightViewportID      ImGuiID
}

struct ImGuiStackLevelInfo {
	iD              ImGuiID
	queryFrameCount ImS8
	querySuccess    bool
	dataType        ImGuiDataType
	desc            [57]i8
}

struct ImVector_ImGuiStackLevelInfo {
	size     int
	capacity int
	data     &ImGuiStackLevelInfo
}

struct ImGuiContextHookCallback {
	lastActiveFrame         int
	stackLevel              int
	queryId                 ImGuiID
	results                 ImVector_ImGuiStackLevelInfo
	copyToClipboardOnCtrlC  bool
	copyToClipboardLastTime f32
	resultPathBuf           ImGuiTextBuffer
}

enum ImGuiContextHookType {
	new_frame_pre
	new_frame_post
	end_frame_pre
	end_frame_post
	render_pre
	render_post
	shutdown
	pending_removal_
}

struct ImGuiContextHook {
	hookId   ImGuiID
	type     ImGuiContextHookType
	owner    ImGuiID
	callback ImGuiContextHookCallback
	userData voidptr
}

struct ImVector_ImGuiInputEvent {
	size     int
	capacity int
	data     &C.ImGuiInputEvent
}

struct ImVector_ImGuiWindowStackData {
	size     int
	capacity int
	data     &ImGuiWindowStackData
}

struct ImVector_ImGuiColorMod {
	size     int
	capacity int
	data     &ImGuiColorMod
}

struct ImVector_ImGuiStyleMod {
	size     int
	capacity int
	data     &ImGuiStyleMod
}

struct ImVector_ImGuiFocusScopeData {
	size     int
	capacity int
	data     &ImGuiFocusScopeData
}

struct ImVector_ImGuiItemFlags {
	size     int
	capacity int
	data     &ImGuiItemFlags
}

struct ImVector_ImGuiGroupData {
	size     int
	capacity int
	data     &ImGuiGroupData
}

struct ImVector_ImGuiPopupData {
	size     int
	capacity int
	data     &ImGuiPopupData
}

struct ImVector_ImGuiTreeNodeStackData {
	size     int
	capacity int
	data     &ImGuiTreeNodeStackData
}

struct ImVector_ImGuiViewportPPtr {
	size     int
	capacity int
	data     &&ImGuiViewportP
}

struct ImVector_unsigned_char {
	size     int
	capacity int
	data     &u8
}

struct ImVector_ImGuiListClipperData {
	size     int
	capacity int
	data     &ImGuiListClipperData
}

struct ImVector_ImGuiTableTempData {
	size     int
	capacity int
	data     &ImGuiTableTempData
}

struct ImVector_ImGuiTable {
	size     int
	capacity int
	data     &ImGuiTable
}

struct ImPool_ImGuiTable {
	buf        ImVector_ImGuiTable
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImGuiTabBar {
	size     int
	capacity int
	data     &C.ImGuiTabBar
}

struct ImPool_ImGuiTabBar {
	buf        ImVector_ImGuiTabBar
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImGuiPtrOrIndex {
	size     int
	capacity int
	data     &ImGuiPtrOrIndex
}

struct ImVector_ImGuiShrinkWidthItem {
	size     int
	capacity int
	data     &ImGuiShrinkWidthItem
}

struct ImVector_ImGuiMultiSelectTempData {
	size     int
	capacity int
	data     &ImGuiMultiSelectTempData
}

struct ImVector_ImGuiMultiSelectState {
	size     int
	capacity int
	data     &ImGuiMultiSelectState
}

struct ImPool_ImGuiMultiSelectState {
	buf        ImVector_ImGuiMultiSelectState
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImGuiID {
	size     int
	capacity int
	data     &ImGuiID
}

struct ImVector_ImGuiSettingsHandler {
	size     int
	capacity int
	data     &ImGuiSettingsHandler
}

struct ImChunkStream_ImGuiWindowSettings {
	buf ImVector_char
}

struct ImChunkStream_ImGuiTableSettings {
	buf ImVector_char
}

struct ImVector_ImGuiContextHook {
	size     int
	capacity int
	data     &ImGuiContextHook
}

struct ImGuiContext {
	initialized                        bool
	fontAtlasOwnedByContext            bool
	iO                                 ImGuiIO
	platformIO                         ImGuiPlatformIO
	style                              ImGuiStyle
	configFlagsCurrFrame               ImGuiConfigFlags
	configFlagsLastFrame               ImGuiConfigFlags
	font                               &ImFont
	fontSize                           f32
	fontBaseSize                       f32
	fontScale                          f32
	currentDpiScale                    f32
	drawListSharedData                 ImDrawListSharedData
	time                               f64
	frameCount                         int
	frameCountEnded                    int
	frameCountPlatformEnded            int
	frameCountRendered                 int
	withinEndChildID                   ImGuiID
	withinFrameScope                   bool
	withinFrameScopeWithImplicitWindow bool
	gcCompactAll                       bool
	testEngineHookItems                bool
	testEngine                         voidptr
	contextName                        [16]i8
	inputEventsQueue                   ImVector_ImGuiInputEvent
	inputEventsTrail                   ImVector_ImGuiInputEvent
	inputEventsNextMouseSource         ImGuiMouseSource
	inputEventsNextEventId             ImU32
	windows                            ImVector_ImGuiWindowPtr
	windowsFocusOrder                  ImVector_ImGuiWindowPtr
	windowsTempSortBuffer              ImVector_ImGuiWindowPtr
	currentWindowStack                 ImVector_ImGuiWindowStackData
	windowsById                        ImGuiStorage
	windowsActiveCount                 int
	windowsBorderHoverPadding          f32
	debugBreakInWindow                 ImGuiID
	currentWindow                      &ImGuiWindow
	hoveredWindow                      &ImGuiWindow
	hoveredWindowUnderMovingWindow     &ImGuiWindow
	hoveredWindowBeforeClear           &ImGuiWindow
	movingWindow                       &ImGuiWindow
	wheelingWindow                     &ImGuiWindow
	wheelingWindowRefMousePos          ImVec2
	wheelingWindowStartFrame           int
	wheelingWindowScrolledFrame        int
	wheelingWindowReleaseTimer         f32
	wheelingWindowWheelRemainder       ImVec2
	wheelingAxisAvg                    ImVec2
	debugDrawIdConflicts               ImGuiID
	debugHookIdInfo                    ImGuiID
	hoveredId                          ImGuiID
	hoveredIdPreviousFrame             ImGuiID
	hoveredIdPreviousFrameItemCount    int
	hoveredIdTimer                     f32
	hoveredIdNotActiveTimer            f32
	hoveredIdAllowOverlap              bool
	hoveredIdIsDisabled                bool
	itemUnclipByLog                    bool
	activeId                           ImGuiID
	activeIdIsAlive                    ImGuiID
	activeIdTimer                      f32
	activeIdIsJustActivated            bool
	activeIdAllowOverlap               bool
	activeIdNoClearOnFocusLoss         bool
	activeIdHasBeenPressedBefore       bool
	activeIdHasBeenEditedBefore        bool
	activeIdHasBeenEditedThisFrame     bool
	activeIdFromShortcut               bool
	activeIdMouseButton                int
	activeIdClickOffset                ImVec2
	activeIdWindow                     &ImGuiWindow
	activeIdSource                     ImGuiInputSource
	activeIdPreviousFrame              ImGuiID
	deactivatedItemData                ImGuiDeactivatedItemData
	activeIdValueOnActivation          ImGuiDataTypeStorage
	lastActiveId                       ImGuiID
	lastActiveIdTimer                  f32
	lastKeyModsChangeTime              f64
	lastKeyModsChangeFromNoneTime      f64
	lastKeyboardKeyPressTime           f64
	keysMayBeCharInput                 ImBitArrayForNamedKeys
	keysOwnerData                      [155]ImGuiKeyOwnerData
	keysRoutingTable                   ImGuiKeyRoutingTable
	activeIdUsingNavDirMask            ImU32
	activeIdUsingAllKeyboardKeys       bool
	debugBreakInShortcutRouting        ImGuiKeyChord
	currentFocusScopeId                ImGuiID
	currentItemFlags                   ImGuiItemFlags
	debugLocateId                      ImGuiID
	nextItemData                       ImGuiNextItemData
	lastItemData                       ImGuiLastItemData
	nextWindowData                     ImGuiNextWindowData
	debugShowGroupRects                bool
	debugFlashStyleColorIdx            ImGuiCol
	colorStack                         ImVector_ImGuiColorMod
	styleVarStack                      ImVector_ImGuiStyleMod
	fontStack                          ImVector_ImFontPtr
	focusScopeStack                    ImVector_ImGuiFocusScopeData
	itemFlagsStack                     ImVector_ImGuiItemFlags
	groupStack                         ImVector_ImGuiGroupData
	openPopupStack                     ImVector_ImGuiPopupData
	beginPopupStack                    ImVector_ImGuiPopupData
	treeNodeStack                      ImVector_ImGuiTreeNodeStackData
	viewports                          ImVector_ImGuiViewportPPtr
	currentViewport                    &ImGuiViewportP
	mouseViewport                      &ImGuiViewportP
	mouseLastHoveredViewport           &ImGuiViewportP
	platformLastFocusedViewportId      ImGuiID
	fallbackMonitor                    ImGuiPlatformMonitor
	platformMonitorsFullWorkRect       C.ImRect
	viewportCreatedCount               int
	platformWindowsCreatedCount        int
	viewportFocusedStampCount          int
	navCursorVisible                   bool
	navHighlightItemUnderNav           bool
	navMousePosDirty                   bool
	navIdIsAlive                       bool
	navId                              ImGuiID
	navWindow                          &ImGuiWindow
	navFocusScopeId                    ImGuiID
	navLayer                           ImGuiNavLayer
	navActivateId                      ImGuiID
	navActivateDownId                  ImGuiID
	navActivatePressedId               ImGuiID
	navActivateFlags                   ImGuiActivateFlags
	navFocusRoute                      ImVector_ImGuiFocusScopeData
	navHighlightActivatedId            ImGuiID
	navHighlightActivatedTimer         f32
	navNextActivateId                  ImGuiID
	navNextActivateFlags               ImGuiActivateFlags
	navInputSource                     ImGuiInputSource
	navLastValidSelectionUserData      ImGuiSelectionUserData
	navCursorHideFrames                ImS8
	navAnyRequest                      bool
	navInitRequest                     bool
	navInitRequestFromMove             bool
	navInitResult                      ImGuiNavItemData
	navMoveSubmitted                   bool
	navMoveScoringItems                bool
	navMoveForwardToNextFrame          bool
	navMoveFlags                       ImGuiNavMoveFlags
	navMoveScrollFlags                 ImGuiScrollFlags
	navMoveKeyMods                     ImGuiKeyChord
	navMoveDir                         ImGuiDir
	navMoveDirForDebug                 ImGuiDir
	navMoveClipDir                     ImGuiDir
	navScoringRect                     C.ImRect
	navScoringNoClipRect               C.ImRect
	navScoringDebugCount               int
	navTabbingDir                      int
	navTabbingCounter                  int
	navMoveResultLocal                 ImGuiNavItemData
	navMoveResultLocalVisible          ImGuiNavItemData
	navMoveResultOther                 ImGuiNavItemData
	navTabbingResultFirst              ImGuiNavItemData
	navJustMovedFromFocusScopeId       ImGuiID
	navJustMovedToId                   ImGuiID
	navJustMovedToFocusScopeId         ImGuiID
	navJustMovedToKeyMods              ImGuiKeyChord
	navJustMovedToIsTabbing            bool
	navJustMovedToHasSelectionData     bool
	configNavWindowingKeyNext          ImGuiKeyChord
	configNavWindowingKeyPrev          ImGuiKeyChord
	navWindowingTarget                 &ImGuiWindow
	navWindowingTargetAnim             &ImGuiWindow
	navWindowingListWindow             &ImGuiWindow
	navWindowingTimer                  f32
	navWindowingHighlightAlpha         f32
	navWindowingToggleLayer            bool
	navWindowingToggleKey              ImGuiKey
	navWindowingAccumDeltaPos          ImVec2
	navWindowingAccumDeltaSize         ImVec2
	dimBgRatio                         f32
	dragDropActive                     bool
	dragDropWithinSource               bool
	dragDropWithinTarget               bool
	dragDropSourceFlags                ImGuiDragDropFlags
	dragDropSourceFrameCount           int
	dragDropMouseButton                int
	dragDropPayload                    ImGuiPayload
	dragDropTargetRect                 C.ImRect
	dragDropTargetClipRect             C.ImRect
	dragDropTargetId                   ImGuiID
	dragDropAcceptFlags                ImGuiDragDropFlags
	dragDropAcceptIdCurrRectSurface    f32
	dragDropAcceptIdCurr               ImGuiID
	dragDropAcceptIdPrev               ImGuiID
	dragDropAcceptFrameCount           int
	dragDropHoldJustPressedId          ImGuiID
	dragDropPayloadBufHeap             ImVector_unsigned_char
	dragDropPayloadBufLocal            [16]u8
	clipperTempDataStacked             int
	clipperTempData                    ImVector_ImGuiListClipperData
	currentTable                       &ImGuiTable
	debugBreakInTable                  ImGuiID
	tablesTempDataStacked              int
	tablesTempData                     ImVector_ImGuiTableTempData
	tables                             ImPool_ImGuiTable
	tablesLastTimeActive               ImVector_float
	drawChannelsTempMergeBuffer        ImVector_ImDrawChannel
	currentTabBar                      &C.ImGuiTabBar
	tabBars                            ImPool_ImGuiTabBar
	currentTabBarStack                 ImVector_ImGuiPtrOrIndex
	shrinkWidthBuffer                  ImVector_ImGuiShrinkWidthItem
	boxSelectState                     ImGuiBoxSelectState
	currentMultiSelect                 &ImGuiMultiSelectTempData
	multiSelectTempDataStacked         int
	multiSelectTempData                ImVector_ImGuiMultiSelectTempData
	multiSelectStorage                 ImPool_ImGuiMultiSelectState
	hoverItemDelayId                   ImGuiID
	hoverItemDelayIdPreviousFrame      ImGuiID
	hoverItemDelayTimer                f32
	hoverItemDelayClearTimer           f32
	hoverItemUnlockedStationaryId      ImGuiID
	hoverWindowUnlockedStationaryId    ImGuiID
	mouseCursor                        ImGuiMouseCursor
	mouseStationaryTimer               f32
	mouseLastValidPos                  ImVec2
	inputTextState                     ImGuiInputTextState
	inputTextDeactivatedState          ImGuiInputTextDeactivatedState
	inputTextPasswordFont              ImFont
	tempInputId                        ImGuiID
	dataTypeZeroValue                  ImGuiDataTypeStorage
	beginMenuDepth                     int
	beginComboDepth                    int
	colorEditOptions                   ImGuiColorEditFlags
	colorEditCurrentID                 ImGuiID
	colorEditSavedID                   ImGuiID
	colorEditSavedHue                  f32
	colorEditSavedSat                  f32
	colorEditSavedColor                ImU32
	colorPickerRef                     C.ImVec4
	comboPreviewData                   ImGuiComboPreviewData
	windowResizeBorderExpectedRect     C.ImRect
	windowResizeRelativeMode           bool
	scrollbarSeekMode                  i16
	scrollbarClickDeltaToGrabCenter    f32
	sliderGrabClickOffset              f32
	sliderCurrentAccum                 f32
	sliderCurrentAccumDirty            bool
	dragCurrentAccumDirty              bool
	dragCurrentAccum                   f32
	dragSpeedDefaultRatio              f32
	disabledAlphaBackup                f32
	disabledStackSize                  i16
	tooltipOverrideCount               i16
	tooltipPreviousWindow              &ImGuiWindow
	clipboardHandlerData               ImVector_char
	menusIdSubmittedThisFrame          ImVector_ImGuiID
	typingSelectState                  ImGuiTypingSelectState
	platformImeData                    ImGuiPlatformImeData
	platformImeDataPrev                ImGuiPlatformImeData
	platformImeViewport                ImGuiID
	dockContext                        ImGuiDockContext
	dockNodeWindowMenuHandler          fn (&ImGuiContext, &ImGuiDockNode, &C.ImGuiTabBar)
	settingsLoaded                     bool
	settingsDirtyTimer                 f32
	settingsIniData                    ImGuiTextBuffer
	settingsHandlers                   ImVector_ImGuiSettingsHandler
	settingsWindows                    ImChunkStream_ImGuiWindowSettings
	settingsTables                     ImChunkStream_ImGuiTableSettings
	hooks                              ImVector_ImGuiContextHook
	hookIdNext                         ImGuiID
	localizationTable                  [13]&i8
	logEnabled                         bool
	logFlags                           ImGuiLogFlags
	logWindow                          &ImGuiWindow
	logFile                            ImFileHandle
	logBuffer                          ImGuiTextBuffer
	logNextPrefix                      &i8
	logNextSuffix                      &i8
	logLinePosY                        f32
	logLineFirstItem                   bool
	logDepthRef                        int
	logDepthToExpand                   int
	logDepthToExpandDefault            int
	errorCallback                      ImGuiErrorCallback
	errorCallbackUserData              voidptr
	errorTooltipLockedPos              ImVec2
	errorFirst                         bool
	errorCountCurrentFrame             int
	stackSizesInNewFrame               ImGuiErrorRecoveryState
	stackSizesInBeginForCurrentWindow  &ImGuiErrorRecoveryState
	debugDrawIdConflictsCount          int
	debugLogFlags                      ImGuiDebugLogFlags
	debugLogBuf                        ImGuiTextBuffer
	debugLogIndex                      ImGuiTextIndex
	debugLogSkippedErrors              int
	debugLogAutoDisableFlags           ImGuiDebugLogFlags
	debugLogAutoDisableFrames          ImU8
	debugLocateFrames                  ImU8
	debugBreakInLocateId               bool
	debugBreakKeyChord                 ImGuiKeyChord
	debugBeginReturnValueCullDepth     ImS8
	debugItemPickerActive              bool
	debugItemPickerMouseButton         ImU8
	debugItemPickerBreakId             ImGuiID
	debugFlashStyleColorTime           f32
	debugFlashStyleColorBackup         C.ImVec4
	debugMetricsConfig                 ImGuiMetricsConfig
	debugIDStackTool                   C.ImGuiIDStackTool
	debugAllocInfo                     ImGuiDebugAllocInfo
	debugHoveredDockNode               &ImGuiDockNode
	framerateSecPerFrame               [60]f32
	framerateSecPerFrameIdx            int
	framerateSecPerFrameCount          int
	framerateSecPerFrameAccum          f32
	wantCaptureMouseNextFrame          int
	wantCaptureKeyboardNextFrame       int
	wantTextInputNextFrame             int
	tempBuffer                         ImVector_char
	tempKeychordName                   [64]i8
}

struct ImGuiWindowTempData {
	cursorPos                 ImVec2
	cursorPosPrevLine         ImVec2
	cursorStartPos            ImVec2
	cursorMaxPos              ImVec2
	idealMaxPos               ImVec2
	currLineSize              ImVec2
	prevLineSize              ImVec2
	currLineTextBaseOffset    f32
	prevLineTextBaseOffset    f32
	isSameLine                bool
	isSetPos                  bool
	indent                    ImVec1
	columnsOffset             ImVec1
	groupOffset               ImVec1
	cursorStartPosLossyness   ImVec2
	navLayerCurrent           ImGuiNavLayer
	navLayersActiveMask       i16
	navLayersActiveMaskNext   i16
	navIsScrollPushableX      bool
	navHideHighlightOneFrame  bool
	navWindowHasScrollY       bool
	menuBarAppending          bool
	menuBarOffset             ImVec2
	menuColumns               ImGuiMenuColumns
	treeDepth                 int
	treeHasStackDataDepthMask ImU32
	childWindows              ImVector_ImGuiWindowPtr
	stateStorage              &ImGuiStorage
	currentColumns            &ImGuiOldColumns
	currentTableIdx           int
	layoutType                ImGuiLayoutType
	parentLayoutType          ImGuiLayoutType
	modalDimBgColor           ImU32
	windowItemStatusFlags     ImGuiItemStatusFlags
	childItemStatusFlags      ImGuiItemStatusFlags
	dockTabItemStatusFlags    ImGuiItemStatusFlags
	dockTabItemRect           C.ImRect
	itemWidth                 f32
	textWrapPos               f32
	itemWidthStack            ImVector_float
	textWrapPosStack          ImVector_float
}

struct ImVector_ImGuiOldColumns {
	size     int
	capacity int
	data     &ImGuiOldColumns
}

struct ImGuiWindow {
	ctx                                &ImGuiContext
	name                               &i8
	iD                                 ImGuiID
	flags                              ImGuiWindowFlags
	flagsPreviousFrame                 ImGuiWindowFlags
	childFlags                         ImGuiChildFlags
	windowClass                        ImGuiWindowClass
	viewport                           &ImGuiViewportP
	viewportId                         ImGuiID
	viewportPos                        ImVec2
	viewportAllowPlatformMonitorExtend int
	pos                                ImVec2
	size                               ImVec2
	sizeFull                           ImVec2
	contentSize                        ImVec2
	contentSizeIdeal                   ImVec2
	contentSizeExplicit                ImVec2
	windowPadding                      ImVec2
	windowRounding                     f32
	windowBorderSize                   f32
	titleBarHeight                     f32
	menuBarHeight                      f32
	decoOuterSizeX1                    f32
	decoOuterSizeY1                    f32
	decoOuterSizeX2                    f32
	decoOuterSizeY2                    f32
	decoInnerSizeX1                    f32
	decoInnerSizeY1                    f32
	nameBufLen                         int
	moveId                             ImGuiID
	tabId                              ImGuiID
	childId                            ImGuiID
	popupId                            ImGuiID
	scroll                             ImVec2
	scrollMax                          ImVec2
	scrollTarget                       ImVec2
	scrollTargetCenterRatio            ImVec2
	scrollTargetEdgeSnapDist           ImVec2
	scrollbarSizes                     ImVec2
	scrollbarX                         bool
	scrollbarY                         bool
	scrollbarXStabilizeEnabled         bool
	scrollbarXStabilizeToggledHistory  ImU8
	viewportOwned                      bool
	active                             bool
	wasActive                          bool
	writeAccessed                      bool
	collapsed                          bool
	wantCollapseToggle                 bool
	skipItems                          bool
	skipRefresh                        bool
	appearing                          bool
	hidden                             bool
	isFallbackWindow                   bool
	isExplicitChild                    bool
	hasCloseButton                     bool
	resizeBorderHovered                i8
	resizeBorderHeld                   i8
	beginCount                         i16
	beginCountPreviousFrame            i16
	beginOrderWithinParent             i16
	beginOrderWithinContext            i16
	focusOrder                         i16
	autoFitFramesX                     ImS8
	autoFitFramesY                     ImS8
	autoFitOnlyGrows                   bool
	autoPosLastDirection               ImGuiDir
	hiddenFramesCanSkipItems           ImS8
	hiddenFramesCannotSkipItems        ImS8
	hiddenFramesForRenderOnly          ImS8
	disableInputsFrames                ImS8
	setWindowPosAllowFlags             ImGuiCond
	setWindowSizeAllowFlags            ImGuiCond
	setWindowCollapsedAllowFlags       ImGuiCond
	setWindowDockAllowFlags            ImGuiCond
	setWindowPosVal                    ImVec2
	setWindowPosPivot                  ImVec2
	iDStack                            ImVector_ImGuiID
	dC                                 ImGuiWindowTempData
	outerRectClipped                   C.ImRect
	innerRect                          C.ImRect
	innerClipRect                      C.ImRect
	workRect                           C.ImRect
	parentWorkRect                     C.ImRect
	clipRect                           C.ImRect
	contentRegionRect                  C.ImRect
	hitTestHoleSize                    ImVec2ih
	hitTestHoleOffset                  ImVec2ih
	lastFrameActive                    int
	lastFrameJustFocused               int
	lastTimeActive                     f32
	itemWidthDefault                   f32
	stateStorage                       ImGuiStorage
	columnsStorage                     ImVector_ImGuiOldColumns
	fontWindowScale                    f32
	fontWindowScaleParents             f32
	fontDpiScale                       f32
	fontRefSize                        f32
	settingsOffset                     int
	drawList                           &ImDrawList
	drawListInst                       ImDrawList
	parentWindow                       &ImGuiWindow
	parentWindowInBeginStack           &ImGuiWindow
	rootWindow                         &ImGuiWindow
	rootWindowPopupTree                &ImGuiWindow
	rootWindowDockTree                 &ImGuiWindow
	rootWindowForTitleBarHighlight     &ImGuiWindow
	rootWindowForNav                   &ImGuiWindow
	parentWindowForFocusRoute          &ImGuiWindow
	navLastChildNavWindow              &ImGuiWindow
	navLastIds                         [2]ImGuiID
	navRectRel                         [2]C.ImRect
	navPreferredScoringPosRel          [2]ImVec2
	navRootFocusScopeId                ImGuiID
	memoryDrawListIdxCapacity          int
	memoryDrawListVtxCapacity          int
	memoryCompacted                    bool
	dockIsActive                       bool
	dockNodeIsVisible                  bool
	dockTabIsVisible                   bool
	dockTabWantClose                   bool
	dockOrder                          i16
	dockStyle                          ImGuiWindowDockStyle
	dockNode                           &ImGuiDockNode
	dockNodeAsHost                     &ImGuiDockNode
	dockId                             ImGuiID
}

enum ImGuiTabBarFlagsPrivate_ {
	dock_node     = 1 << 20
	is_focused    = 1 << 21
	save_settings = 1 << 22
}

enum ImGuiTabItemFlagsPrivate_ {
	section_mask_   = 1 << 6 | 1 << 7
	no_close_button = 1 << 20
	button          = 1 << 21
	invisible       = 1 << 22
	unsorted        = 1 << 23
}

struct ImGuiTabItem {
	iD                ImGuiID
	flags             ImGuiTabItemFlags
	window            &ImGuiWindow
	lastFrameVisible  int
	lastFrameSelected int
	offset            f32
	width             f32
	contentWidth      f32
	requestedWidth    f32
	nameOffset        ImS32
	beginOrder        ImS16
	indexDuringLayout ImS16
	wantClose         bool
}

struct ImVector_ImGuiTabItem {
	size     int
	capacity int
	data     &ImGuiTabItem
}

struct ImGuiTableColumnIdx {
	window                          &ImGuiWindow
	tabs                            ImVector_ImGuiTabItem
	flags                           ImGuiTabBarFlags
	iD                              ImGuiID
	selectedTabId                   ImGuiID
	nextSelectedTabId               ImGuiID
	visibleTabId                    ImGuiID
	currFrameVisible                int
	prevFrameVisible                int
	barRect                         C.ImRect
	currTabsContentsHeight          f32
	prevTabsContentsHeight          f32
	widthAllTabs                    f32
	widthAllTabsIdeal               f32
	scrollingAnim                   f32
	scrollingTarget                 f32
	scrollingTargetDistToVisibility f32
	scrollingSpeed                  f32
	scrollingRectMinX               f32
	scrollingRectMaxX               f32
	separatorMinX                   f32
	separatorMaxX                   f32
	reorderRequestTabId             ImGuiID
	reorderRequestOffset            ImS16
	beginCount                      ImS8
	wantLayout                      bool
	visibleTabWasSubmitted          bool
	tabsAddedNew                    bool
	tabsActiveCount                 ImS16
	lastTabItemIdx                  ImS16
	itemSpacingY                    f32
	framePadding                    ImVec2
	backupCursorPos                 ImVec2
	tabsNames                       ImGuiTextBuffer
}

type ImGuiTableDrawChannelIdx = u16

struct ImGuiTableColumn {
	flags                    ImGuiTableColumnFlags
	widthGiven               f32
	minX                     f32
	maxX                     f32
	widthRequest             f32
	widthAuto                f32
	widthMax                 f32
	stretchWeight            f32
	initStretchWeightOrWidth f32
	clipRect                 C.ImRect
	userID                   ImGuiID
	workMinX                 f32
	workMaxX                 f32
	itemWidth                f32
	contentMaxXFrozen        f32
	contentMaxXUnfrozen      f32
	contentMaxXHeadersUsed   f32
	contentMaxXHeadersIdeal  f32
	nameOffset               ImS16
	displayOrder             ImGuiTableColumnIdx
	indexWithinEnabledSet    ImGuiTableColumnIdx
	prevEnabledColumn        ImGuiTableColumnIdx
	nextEnabledColumn        ImGuiTableColumnIdx
	sortOrder                ImGuiTableColumnIdx
	drawChannelCurrent       ImGuiTableDrawChannelIdx
	drawChannelFrozen        ImGuiTableDrawChannelIdx
	drawChannelUnfrozen      ImGuiTableDrawChannelIdx
	isEnabled                bool
	isUserEnabled            bool
	isUserEnabledNextFrame   bool
	isVisibleX               bool
	isVisibleY               bool
	isRequestOutput          bool
	isSkipItems              bool
	isPreserveWidthAuto      bool
	navLayerCurrent          ImS8
	autoFitQueue             ImU8
	cannotSkipItemsQueue     ImU8
	sortDirection            ImU8
	sortDirectionsAvailCount ImU8
	sortDirectionsAvailMask  ImU8
	sortDirectionsAvailList  ImU8
}

struct ImGuiTableCellData {
	bgColor ImU32
	column  ImGuiTableColumnIdx
}

struct ImGuiTableHeaderData {
	index     ImGuiTableColumnIdx
	textColor ImU32
	bgColor0  ImU32
	bgColor1  ImU32
}

struct ImGuiTableInstanceData {
	tableInstanceID         ImGuiID
	lastOuterHeight         f32
	lastTopHeadersRowHeight f32
	lastFrozenHeight        f32
	hoveredRowLast          int
	hoveredRowNext          int
}

struct ImSpan_ImGuiTableColumn {
	data    &ImGuiTableColumn
	dataEnd &ImGuiTableColumn
}

struct ImSpan_ImGuiTableColumnIdx {
	data    &ImGuiTableColumnIdx
	dataEnd &ImGuiTableColumnIdx
}

struct ImSpan_ImGuiTableCellData {
	data    &ImGuiTableCellData
	dataEnd &ImGuiTableCellData
}

struct ImVector_ImGuiTableInstanceData {
	size     int
	capacity int
	data     &ImGuiTableInstanceData
}

struct ImVector_ImGuiTableColumnSortSpecs {
	size     int
	capacity int
	data     &ImGuiTableColumnSortSpecs
}

struct ImGuiTable {
	iD                         ImGuiID
	flags                      ImGuiTableFlags
	rawData                    voidptr
	tempData                   &ImGuiTableTempData
	columns                    ImSpan_ImGuiTableColumn
	displayOrderToIndex        ImSpan_ImGuiTableColumnIdx
	rowCellData                ImSpan_ImGuiTableCellData
	enabledMaskByDisplayOrder  ImBitArrayPtr
	enabledMaskByIndex         ImBitArrayPtr
	visibleMaskByIndex         ImBitArrayPtr
	settingsLoadedFlags        ImGuiTableFlags
	settingsOffset             int
	lastFrameActive            int
	columnsCount               int
	currentRow                 int
	currentColumn              int
	instanceCurrent            ImS16
	instanceInteracted         ImS16
	rowPosY1                   f32
	rowPosY2                   f32
	rowMinHeight               f32
	rowCellPaddingY            f32
	rowTextBaseline            f32
	rowIndentOffsetX           f32
	rowFlags                   ImGuiTableRowFlags
	lastRowFlags               ImGuiTableRowFlags
	rowBgColorCounter          int
	rowBgColor                 [2]ImU32
	borderColorStrong          ImU32
	borderColorLight           ImU32
	borderX1                   f32
	borderX2                   f32
	hostIndentX                f32
	minColumnWidth             f32
	outerPaddingX              f32
	cellPaddingX               f32
	cellSpacingX1              f32
	cellSpacingX2              f32
	innerWidth                 f32
	columnsGivenWidth          f32
	columnsAutoFitWidth        f32
	columnsStretchSumWeights   f32
	resizedColumnNextWidth     f32
	resizeLockMinContentsX2    f32
	refScale                   f32
	angledHeadersHeight        f32
	angledHeadersSlope         f32
	outerRect                  C.ImRect
	innerRect                  C.ImRect
	workRect                   C.ImRect
	innerClipRect              C.ImRect
	bgClipRect                 C.ImRect
	bg0ClipRectForDrawCmd      C.ImRect
	bg2ClipRectForDrawCmd      C.ImRect
	hostClipRect               C.ImRect
	hostBackupInnerClipRect    C.ImRect
	outerWindow                &ImGuiWindow
	innerWindow                &ImGuiWindow
	columnsNames               ImGuiTextBuffer
	drawSplitter               &ImDrawListSplitter
	instanceDataFirst          ImGuiTableInstanceData
	instanceDataExtra          ImVector_ImGuiTableInstanceData
	sortSpecsSingle            ImGuiTableColumnSortSpecs
	sortSpecsMulti             ImVector_ImGuiTableColumnSortSpecs
	sortSpecs                  ImGuiTableSortSpecs
	sortSpecsCount             ImGuiTableColumnIdx
	columnsEnabledCount        ImGuiTableColumnIdx
	columnsEnabledFixedCount   ImGuiTableColumnIdx
	declColumnsCount           ImGuiTableColumnIdx
	angledHeadersCount         ImGuiTableColumnIdx
	hoveredColumnBody          ImGuiTableColumnIdx
	hoveredColumnBorder        ImGuiTableColumnIdx
	highlightColumnHeader      ImGuiTableColumnIdx
	autoFitSingleColumn        ImGuiTableColumnIdx
	resizedColumn              ImGuiTableColumnIdx
	lastResizedColumn          ImGuiTableColumnIdx
	heldHeaderColumn           ImGuiTableColumnIdx
	reorderColumn              ImGuiTableColumnIdx
	reorderColumnDir           ImGuiTableColumnIdx
	leftMostEnabledColumn      ImGuiTableColumnIdx
	rightMostEnabledColumn     ImGuiTableColumnIdx
	leftMostStretchedColumn    ImGuiTableColumnIdx
	rightMostStretchedColumn   ImGuiTableColumnIdx
	contextPopupColumn         ImGuiTableColumnIdx
	freezeRowsRequest          ImGuiTableColumnIdx
	freezeRowsCount            ImGuiTableColumnIdx
	freezeColumnsRequest       ImGuiTableColumnIdx
	freezeColumnsCount         ImGuiTableColumnIdx
	rowCellDataCurrent         ImGuiTableColumnIdx
	dummyDrawChannel           ImGuiTableDrawChannelIdx
	bg2DrawChannelCurrent      ImGuiTableDrawChannelIdx
	bg2DrawChannelUnfrozen     ImGuiTableDrawChannelIdx
	navLayer                   ImS8
	isLayoutLocked             bool
	isInsideRow                bool
	isInitializing             bool
	isSortSpecsDirty           bool
	isUsingHeaders             bool
	isContextPopupOpen         bool
	disableDefaultContextMenu  bool
	isSettingsRequestLoad      bool
	isSettingsDirty            bool
	isDefaultDisplayOrder      bool
	isResetAllRequest          bool
	isResetDisplayOrderRequest bool
	isUnfrozenRows             bool
	isDefaultSizingPolicy      bool
	isActiveIdAliveBeforeTable bool
	isActiveIdInTable          bool
	hasScrollbarYCurr          bool
	hasScrollbarYPrev          bool
	memoryCompacted            bool
	hostSkipItems              bool
}

struct ImVector_ImGuiTableHeaderData {
	size     int
	capacity int
	data     &ImGuiTableHeaderData
}

struct ImGuiTableTempData {
	tableIndex                   int
	lastTimeActive               f32
	angledHeadersExtraWidth      f32
	angledHeadersRequests        ImVector_ImGuiTableHeaderData
	userOuterSize                ImVec2
	drawSplitter                 ImDrawListSplitter
	hostBackupWorkRect           C.ImRect
	hostBackupParentWorkRect     C.ImRect
	hostBackupPrevLineSize       ImVec2
	hostBackupCurrLineSize       ImVec2
	hostBackupCursorMaxPos       ImVec2
	hostBackupColumnsOffset      ImVec1
	hostBackupItemWidth          f32
	hostBackupItemWidthStackSize int
}

struct ImGuiTableColumnSettings {
	widthOrWeight f32
	userID        ImGuiID
	index         ImGuiTableColumnIdx
	displayOrder  ImGuiTableColumnIdx
	sortOrder     ImGuiTableColumnIdx
	sortDirection ImU8
	isEnabled     ImS8
	isStretch     ImU8
}

struct ImGuiTableSettings {
	iD              ImGuiID
	saveFlags       ImGuiTableFlags
	refScale        f32
	columnsCount    ImGuiTableColumnIdx
	columnsCountMax ImGuiTableColumnIdx
	wantApply       bool
}

struct ImFontBuilderIO {
	fontBuilder_Build fn (&ImFontAtlas) bool
}

// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
/////////////////////////hand written functions
// no LogTextV
// no appendfV
// for getting FLT_MAX in bindings
// for getting FLT_MIN in bindings
// CIMGUI_INCLUDED
// This file is automatically generated by int(generator.lua) from https://int(github.com)/cimgui/cimplot
// based on int(implot.h) file version int(0.17) from implot https://int(github.com)/epezent/implot
// with int(implot_internal.h) api
struct ImVector_ImS16 {
	size     int
	capacity int
	data     &ImS16
}

struct ImVector_ImS32 {
	size     int
	capacity int
	data     &ImS32
}

struct ImVector_ImS64 {
	size     int
	capacity int
	data     &ImS64
}

struct ImVector_ImS8 {
	size     int
	capacity int
	data     &ImS8
}

struct ImVector_ImU64 {
	size     int
	capacity int
	data     &ImU64
}

type ImAxis = int
type Flags = int
type AxisFlags = int
type SubplotFlags = int
type LegendFlags = int
type MouseTextFlags = int
type DragToolFlags = int
type ColormapScaleFlags = int
type ItemFlags = int
type LineFlags = int
type ScatterFlags = int
type StairsFlags = int
type ShadedFlags = int
type BarsFlags = int
type BarGroupsFlags = int
type ErrorBarsFlags = int
type StemsFlags = int
type InfLinesFlags = int
type PieChartFlags = int
type HeatmapFlags = int
type HistogramFlags = int
type DigitalFlags = int
type ImageFlags = int
type TextFlags = int
type DummyFlags = int
type Cond = int
type Col = int
type StyleVar = int
type Scale = int
type Marker = int
type Colormap = int
type Location = int
type Bin = int

enum ImAxis_ {
	x1 = 0
	x2
	x3
	y1
	y2
	y3
	count
}

enum Flags_ {
	none          = 0
	no_title      = 1 << 0
	no_legend     = 1 << 1
	no_mouse_text = 1 << 2
	no_inputs     = 1 << 3
	no_menus      = 1 << 4
	no_box_select = 1 << 5
	no_frame      = 1 << 6
	equal         = 1 << 7
	crosshairs    = 1 << 8
	canvas_only   = 1 << 0 | 1 << 1 | 1 << 4 | 1 << 5 | 1 << 2
}

enum AxisFlags_ {
	none           = 0
	no_label       = 1 << 0
	no_grid_lines  = 1 << 1
	no_tick_marks  = 1 << 2
	no_tick_labels = 1 << 3
	no_initial_fit = 1 << 4
	no_menus       = 1 << 5
	no_side_switch = 1 << 6
	no_highlight   = 1 << 7
	opposite       = 1 << 8
	foreground     = 1 << 9
	invert         = 1 << 10
	auto_fit       = 1 << 11
	range_fit      = 1 << 12
	pan_stretch    = 1 << 13
	lock_min       = 1 << 14
	lock_max       = 1 << 15
	lock           = 1 << 14 | 1 << 15
	no_decorations = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
	aux_default    = 1 << 1 | 1 << 8
}

enum SubplotFlags_ {
	none        = 0
	no_title    = 1 << 0
	no_legend   = 1 << 1
	no_menus    = 1 << 2
	no_resize   = 1 << 3
	no_align    = 1 << 4
	share_items = 1 << 5
	link_rows   = 1 << 6
	link_cols   = 1 << 7
	link_all_x  = 1 << 8
	link_all_y  = 1 << 9
	col_major   = 1 << 10
}

enum LegendFlags_ {
	none              = 0
	no_buttons        = 1 << 0
	no_highlight_item = 1 << 1
	no_highlight_axis = 1 << 2
	no_menus          = 1 << 3
	outside           = 1 << 4
	horizontal        = 1 << 5
	sort              = 1 << 6
}

enum MouseTextFlags_ {
	none        = 0
	no_aux_axes = 1 << 0
	no_format   = 1 << 1
	show_always = 1 << 2
}

enum DragToolFlags_ {
	none       = 0
	no_cursors = 1 << 0
	no_fit     = 1 << 1
	no_inputs  = 1 << 2
	delayed    = 1 << 3
}

enum ColormapScaleFlags_ {
	none     = 0
	no_label = 1 << 0
	opposite = 1 << 1
	invert   = 1 << 2
}

enum ItemFlags_ {
	none      = 0
	no_legend = 1 << 0
	no_fit    = 1 << 1
}

enum LineFlags_ {
	none      = 0
	segments  = 1 << 10
	loop      = 1 << 11
	skip_na_n = 1 << 12
	no_clip   = 1 << 13
	shaded    = 1 << 14
}

enum ScatterFlags_ {
	none    = 0
	no_clip = 1 << 10
}

enum StairsFlags_ {
	none     = 0
	pre_step = 1 << 10
	shaded   = 1 << 11
}

enum ShadedFlags_ {
	none = 0
}

enum BarsFlags_ {
	none       = 0
	horizontal = 1 << 10
}

enum BarGroupsFlags_ {
	none       = 0
	horizontal = 1 << 10
	stacked    = 1 << 11
}

enum ErrorBarsFlags_ {
	none       = 0
	horizontal = 1 << 10
}

enum StemsFlags_ {
	none       = 0
	horizontal = 1 << 10
}

enum InfLinesFlags_ {
	none       = 0
	horizontal = 1 << 10
}

enum PieChartFlags_ {
	none          = 0
	normalize     = 1 << 10
	ignore_hidden = 1 << 11
	exploding     = 1 << 12
}

enum HeatmapFlags_ {
	none      = 0
	col_major = 1 << 10
}

enum HistogramFlags_ {
	none        = 0
	horizontal  = 1 << 10
	cumulative  = 1 << 11
	density     = 1 << 12
	no_outliers = 1 << 13
	col_major   = 1 << 14
}

enum DigitalFlags_ {
	none = 0
}

enum ImageFlags_ {
	none = 0
}

enum TextFlags_ {
	none     = 0
	vertical = 1 << 10
}

enum DummyFlags_ {
	none = 0
}

enum Cond_ {
	none   = 0
	always = 1 << 0
	once   = 1 << 1
}

enum Col_ {
	line
	fill
	marker_outline
	marker_fill
	error_bar
	frame_bg
	plot_bg
	plot_border
	legend_bg
	legend_border
	legend_text
	title_text
	inlay_text
	axis_text
	axis_grid
	axis_tick
	axis_bg
	axis_bg_hovered
	axis_bg_active
	selection
	crosshairs
	count
}

enum StyleVar_ {
	line_weight
	marker
	marker_size
	marker_weight
	fill_alpha
	error_bar_size
	error_bar_weight
	digital_bit_height
	digital_bit_gap
	plot_border_size
	minor_alpha
	major_tick_len
	minor_tick_len
	major_tick_size
	minor_tick_size
	major_grid_size
	minor_grid_size
	plot_padding
	label_padding
	legend_padding
	legend_inner_padding
	legend_spacing
	mouse_pos_padding
	annotation_padding
	fit_padding
	plot_default_size
	plot_min_size
	count
}

enum Scale_ {
	linear = 0
	time
	log10
	sym_log
}

enum Marker_ {
	none = -1
	circle
	square
	diamond
	up
	down
	left
	right
	cross
	plus
	asterisk
	count
}

enum Colormap_ {
	deep     = 0
	dark     = 1
	pastel   = 2
	paired   = 3
	viridis  = 4
	plasma   = 5
	hot      = 6
	cool     = 7
	pink     = 8
	jet      = 9
	twilight = 10
	rd_bu    = 11
	br_bg    = 12
	pi_yg    = 13
	spectral = 14
	greys    = 15
}

enum Location_ {
	center     = 0
	north      = 1 << 0
	south      = 1 << 1
	west       = 1 << 2
	east       = 1 << 3
	north_west = 1 << 0 | 1 << 2
	north_east = 1 << 0 | 1 << 3
	south_west = 1 << 1 | 1 << 2
	south_east = 1 << 1 | 1 << 3
}

enum Bin_ {
	sqrt    = -1
	sturges = -2
	rice    = -3
	scott   = -4
}

struct Point {
	x f64
	y f64
}

struct Range {
	min f64
	max f64
}

struct Rect {
	x Range
	y Range
}

struct Style {
	lineWeight         f32
	marker             int
	markerSize         f32
	markerWeight       f32
	fillAlpha          f32
	errorBarSize       f32
	errorBarWeight     f32
	digitalBitHeight   f32
	digitalBitGap      f32
	plotBorderSize     f32
	minorAlpha         f32
	majorTickLen       ImVec2
	minorTickLen       ImVec2
	majorTickSize      ImVec2
	minorTickSize      ImVec2
	majorGridSize      ImVec2
	minorGridSize      ImVec2
	plotPadding        ImVec2
	labelPadding       ImVec2
	legendPadding      ImVec2
	legendInnerPadding ImVec2
	legendSpacing      ImVec2
	mousePosPadding    ImVec2
	annotationPadding  ImVec2
	fitPadding         ImVec2
	plotDefaultSize    ImVec2
	plotMinSize        ImVec2
	colors             [21]C.ImVec4
	colormap           Colormap
	useLocalTime       bool
	useISO8601         bool
	use24HourClock     bool
}

struct Formatter {
	pan           ImGuiMouseButton
	panMod        int
	fit           ImGuiMouseButton
	select        ImGuiMouseButton
	selectCancel  ImGuiMouseButton
	selectMod     int
	selectHorzMod int
	selectVertMod int
	menu          ImGuiMouseButton
	overrideMod   int
	zoomMod       int
	zoomRate      f32
}

type Getter = fn (int, voidptr) Point

type Transform = fn (f64, voidptr) f64

@[weak]
__global GImPlot &Context

type TimeUnit = int
type DateFmt = int
type TimeFmt = int

enum TimeUnit_ {
	us
	ms
	s
	min
	hr
	day
	mo
	yr
	count
}

enum DateFmt_ {
	none = 0
	day_mo
	day_mo_yr
	mo_yr
	mo
	yr
}

enum TimeFmt_ {
	none = 0
	us
	su_s
	sm_s
	s
	min_sm_s
	hr_min_sm_s
	hr_min_s
	hr_min
	hr
}

type Locator = fn (&Ticker, Range, f32, bool, Formatter, voidptr)

struct DateTimeSpec {
	date           DateFmt
	time           TimeFmt
	useISO8601     bool
	use24HourClock bool
}

struct Time {
	s  C.time_t
	us int
}

struct ImVector_bool {
	size     int
	capacity int
	data     &bool
}

struct ColormapData {
	keys         ImVector_ImU32
	keyCounts    ImVector_int
	keyOffsets   ImVector_int
	tables       ImVector_ImU32
	tableSizes   ImVector_int
	tableOffsets ImVector_int
	text         ImGuiTextBuffer
	textOffsets  ImVector_int
	quals        ImVector_bool
	map          ImGuiStorage
	count        int
}

struct PointError {
	x   f64
	y   f64
	neg f64
	pos f64
}

struct Annotation {
	pos        ImVec2
	offset     ImVec2
	colorBg    ImU32
	colorFg    ImU32
	textOffset int
	clamp      bool
}

struct ImVector_ImPlotAnnotation {
	size     int
	capacity int
	data     &Annotation
}

struct AnnotationCollection {
	annotations ImVector_ImPlotAnnotation
	textBuffer  ImGuiTextBuffer
	size        int
}

struct Tag {
	axis       ImAxis
	value      f64
	colorBg    ImU32
	colorFg    ImU32
	textOffset int
}

struct ImVector_ImPlotTag {
	size     int
	capacity int
	data     &Tag
}

struct TagCollection {
	tags       ImVector_ImPlotTag
	textBuffer ImGuiTextBuffer
	size       int
}

struct Tick {
	plotPos    f64
	pixelPos   f32
	labelSize  ImVec2
	textOffset int
	major      bool
	showLabel  bool
	level      int
	idx        int
}

struct ImVector_ImPlotTick {
	size     int
	capacity int
	data     &Tick
}

struct Ticker {
	ticks      ImVector_ImPlotTick
	textBuffer ImGuiTextBuffer
	maxSize    ImVec2
	lateSize   ImVec2
	levels     int
}

struct Axis {
	iD               ImGuiID
	flags            AxisFlags
	previousFlags    AxisFlags
	range            Range
	rangeCond        Cond
	scale            Scale
	fitExtents       Range
	orthoAxis        &Axis
	constraintRange  Range
	constraintZoom   Range
	ticker           Ticker
	formatter        Formatter
	formatterData    voidptr
	formatSpec       [16]i8
	locator          Locator
	linkedMin        &f64
	linkedMax        &f64
	pickerLevel      int
	pickerTimeMin    Time
	pickerTimeMax    Time
	transformForward Transform
	transformInverse Transform
	transformData    voidptr
	pixelMin         f32
	pixelMax         f32
	scaleMin         f64
	scaleMax         f64
	scaleToPixel     f64
	datum1           f32
	datum2           f32
	hoverRect        C.ImRect
	labelOffset      int
	colorMaj         ImU32
	colorMin         ImU32
	colorTick        ImU32
	colorTxt         ImU32
	colorBg          ImU32
	colorHov         ImU32
	colorAct         ImU32
	colorHiLi        ImU32
	enabled          bool
	vertical         bool
	fitThisFrame     bool
	hasRange         bool
	hasFormatSpec    bool
	showDefaultTicks bool
	hovered          bool
	held             bool
}

struct AlignmentData {
	vertical bool
	padA     f32
	padB     f32
	padAMax  f32
	padBMax  f32
}

struct Item {
	iD              ImGuiID
	color           ImU32
	legendHoverRect C.ImRect
	nameOffset      int
	show            bool
	legendHovered   bool
	seenThisFrame   bool
}

struct Legend {
	flags            LegendFlags
	previousFlags    LegendFlags
	location         Location
	previousLocation Location
	scroll           ImVec2
	indices          ImVector_int
	labels           ImGuiTextBuffer
	rect             C.ImRect
	rectClamped      C.ImRect
	hovered          bool
	held             bool
	canGoInside      bool
}

struct ImVector_ImPlotItem {
	size     int
	capacity int
	data     &Item
}

struct ImPool_ImPlotItem {
	buf        ImVector_ImPlotItem
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ItemGroup {
	iD          ImGuiID
	legend      Legend
	itemPool    ImPool_ImPlotItem
	colormapIdx int
}

struct Plot {
	iD                ImGuiID
	flags             Flags
	previousFlags     Flags
	mouseTextLocation Location
	mouseTextFlags    MouseTextFlags
	axes              [6]Axis
	textBuffer        ImGuiTextBuffer
	items             ItemGroup
	currentX          ImAxis
	currentY          ImAxis
	frameRect         C.ImRect
	canvasRect        C.ImRect
	plotRect          C.ImRect
	axesRect          C.ImRect
	selectRect        C.ImRect
	selectStart       ImVec2
	titleOffset       int
	justCreated       bool
	initialized       bool
	setupLocked       bool
	fitThisFrame      bool
	hovered           bool
	held              bool
	selecting         bool
	selected          bool
	contextLocked     bool
}

struct ImVector_ImPlotAlignmentData {
	size     int
	capacity int
	data     &AlignmentData
}

struct ImVector_ImPlotRange {
	size     int
	capacity int
	data     &Range
}

struct Subplot {
	iD               ImGuiID
	flags            SubplotFlags
	previousFlags    SubplotFlags
	items            ItemGroup
	rows             int
	cols             int
	currentIdx       int
	frameRect        C.ImRect
	gridRect         C.ImRect
	cellSize         ImVec2
	rowAlignmentData ImVector_ImPlotAlignmentData
	colAlignmentData ImVector_ImPlotAlignmentData
	rowRatios        ImVector_float
	colRatios        ImVector_float
	rowLinkData      ImVector_ImPlotRange
	colLinkData      ImVector_ImPlotRange
	tempSizes        [2]f32
	frameHovered     bool
	hasTitle         bool
}

struct NextPlotData {
	rangeCond [6]Cond
	range     [6]Range
	hasRange  [6]bool
	fit       [6]bool
	linkedMin [6]&f64
	linkedMax [6]&f64
}

struct NextItemData {
	colors           [5]C.ImVec4
	lineWeight       f32
	marker           Marker
	markerSize       f32
	markerWeight     f32
	fillAlpha        f32
	errorBarSize     f32
	errorBarWeight   f32
	digitalBitHeight f32
	digitalBitGap    f32
	renderLine       bool
	renderFill       bool
	renderMarkerLine bool
	renderMarkerFill bool
	hasHidden        bool
	hidden           bool
	hiddenCond       Cond
}

struct ImVector_ImPlotPlot {
	size     int
	capacity int
	data     &Plot
}

struct ImPool_ImPlotPlot {
	buf        ImVector_ImPlotPlot
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImPlotSubplot {
	size     int
	capacity int
	data     &Subplot
}

struct ImPool_ImPlotSubplot {
	buf        ImVector_ImPlotSubplot
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImPlotColormap {
	size     int
	capacity int
	data     &Colormap
}

struct ImVector_double {
	size     int
	capacity int
	data     &f64
}

struct ImPool_ImPlotAlignmentData {
	buf        ImVector_ImPlotAlignmentData
	map        ImGuiStorage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct Context {
	plots                 ImPool_ImPlotPlot
	subplots              ImPool_ImPlotSubplot
	currentPlot           &Plot
	currentSubplot        &Subplot
	currentItems          &ItemGroup
	currentItem           &Item
	previousItem          &Item
	cTicker               Ticker
	annotations           AnnotationCollection
	tags                  TagCollection
	style                 Style
	colorModifiers        ImVector_ImGuiColorMod
	styleModifiers        ImVector_ImGuiStyleMod
	colormapData          ColormapData
	colormapModifiers     ImVector_ImPlotColormap
	tm                    C.tm
	tempDouble1           ImVector_double
	tempDouble2           ImVector_double
	tempInt1              ImVector_int
	digitalPlotItemCnt    int
	digitalPlotOffset     int
	nextPlotData          NextPlotData
	nextItemData          NextItemData
	inputMap              InputMap
	openContextThisFrame  bool
	mousePosStringBuilder ImGuiTextBuffer
	sortItems             &ItemGroup
	alignmentData         ImPool_ImPlotAlignmentData
	currentAlignmentH     &AlignmentData
	currentAlignmentV     &AlignmentData
}

struct Point_getter {
	time              Time
	spec              DateTimeSpec
	userFormatter     Formatter
	userFormatterData voidptr
}

// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
// Point getters manually wrapped use this
// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
@[c: 'ImPlotPoint_ImPlotPoint_Nil']
fn point_im_plot_point_nil() &Point

@[c: 'ImPlotPoint_destroy']
fn point_destroy(self &Point)

@[c: 'ImPlotPoint_ImPlotPoint_double']
fn point_im_plot_point_double(_x f64, _y f64) &Point

@[c: 'ImPlotPoint_ImPlotPoint_Vec2']
fn point_im_plot_point_vec2(p ImVec2) &Point

@[c: 'ImPlotRange_ImPlotRange_Nil']
fn range_im_plot_range_nil() &Range

@[c: 'ImPlotRange_destroy']
fn range_destroy(self &Range)

@[c: 'ImPlotRange_ImPlotRange_double']
fn range_im_plot_range_double(_min f64, _max f64) &Range

@[c: 'ImPlotRange_Contains']
fn range_contains(self &Range, value f64) bool

@[c: 'ImPlotRange_Size']
fn range_size(self &Range) f64

@[c: 'ImPlotRange_Clamp']
fn range_clamp(self &Range, value f64) f64

@[c: 'ImPlotRect_ImPlotRect_Nil']
fn rect_im_plot_rect_nil() &Rect

@[c: 'ImPlotRect_destroy']
fn rect_destroy(self &Rect)

@[c: 'ImPlotRect_ImPlotRect_double']
fn rect_im_plot_rect_double(x_min f64, x_max f64, y_min f64, y_max f64) &Rect

@[c: 'ImPlotRect_Contains_PlotPoInt']
fn rect_contains_plot_po_int(self &Rect, p Point) bool

@[c: 'ImPlotRect_Contains_double']
fn rect_contains_double(self &Rect, x f64, y f64) bool

@[c: 'ImPlotRect_Size']
fn rect_size(p_out &Point, self &Rect)

@[c: 'ImPlotRect_Clamp_PlotPoInt']
fn rect_clamp_plot_po_int(p_out &Point, self &Rect, p Point)

@[c: 'ImPlotRect_Clamp_double']
fn rect_clamp_double(p_out &Point, self &Rect, x f64, y f64)

@[c: 'ImPlotRect_Min']
fn rect_min(p_out &Point, self &Rect)

@[c: 'ImPlotRect_Max']
fn rect_max(p_out &Point, self &Rect)

@[c: 'ImPlotStyle_ImPlotStyle']
fn style_im_plot_style() &Style

@[c: 'ImPlotStyle_destroy']
fn style_destroy(self &Style)

@[c: 'ImPlotInputMap_ImPlotInputMap']
fn input_map_im_plot_input_map() &InputMap

@[c: 'ImPlotInputMap_destroy']
fn input_map_destroy(self &InputMap)

@[c: 'ImPlot_CreateContext']
fn create_context() &Context

@[c: 'ImPlot_DestroyContext']
fn destroy_context(ctx &Context)

@[c: 'ImPlot_GetCurrentContext']
fn get_current_context() &Context

@[c: 'ImPlot_SetCurrentContext']
fn set_current_context(ctx &Context)

@[c: 'ImPlot_SetImGuiContext']
fn set_im_gui_context(ctx &ImGuiContext)

@[c: 'ImPlot_BeginPlot']
fn begin_plot(title_id &i8, size ImVec2, flags Flags) bool

@[c: 'ImPlot_EndPlot']
fn end_plot()

@[c: 'ImPlot_BeginSubplots']
fn begin_subplots(title_id &i8, rows int, cols int, size ImVec2, flags SubplotFlags, row_ratios &f32, col_ratios &f32) bool

@[c: 'ImPlot_EndSubplots']
fn end_subplots()

@[c: 'ImPlot_SetupAxis']
fn setup_axis(axis ImAxis, label &i8, flags AxisFlags)

@[c: 'ImPlot_SetupAxisLimits']
fn setup_axis_limits(axis ImAxis, v_min f64, v_max f64, cond Cond)

@[c: 'ImPlot_SetupAxisLinks']
fn setup_axis_links(axis ImAxis, link_min &f64, link_max &f64)

@[c: 'ImPlot_SetupAxisFormat_Str']
fn setup_axis_format_str(axis ImAxis, fmt &i8)

@[c: 'ImPlot_SetupAxisFormat_PlotFormatter']
fn setup_axis_format_plot_formatter(axis ImAxis, formatter Formatter, data voidptr)

@[c: 'ImPlot_SetupAxisTicks_doublePtr']
fn setup_axis_ticks_double_ptr(axis ImAxis, values &f64, n_ticks int, labels &&u8, keep_default bool)

@[c: 'ImPlot_SetupAxisTicks_double']
fn setup_axis_ticks_double(axis ImAxis, v_min f64, v_max f64, n_ticks int, labels &&u8, keep_default bool)

@[c: 'ImPlot_SetupAxisScale_PlotScale']
fn setup_axis_scale_plot_scale(axis ImAxis, scale Scale)

@[c: 'ImPlot_SetupAxisScale_PlotTransform']
fn setup_axis_scale_plot_transform(axis ImAxis, forward Transform, inverse Transform, data voidptr)

@[c: 'ImPlot_SetupAxisLimitsConstraints']
fn setup_axis_limits_constraints(axis ImAxis, v_min f64, v_max f64)

@[c: 'ImPlot_SetupAxisZoomConstraints']
fn setup_axis_zoom_constraints(axis ImAxis, z_min f64, z_max f64)

@[c: 'ImPlot_SetupAxes']
fn setup_axes(x_label &i8, y_label &i8, x_flags AxisFlags, y_flags AxisFlags)

@[c: 'ImPlot_SetupAxesLimits']
fn setup_axes_limits(x_min f64, x_max f64, y_min f64, y_max f64, cond Cond)

@[c: 'ImPlot_SetupLegend']
fn setup_legend(location Location, flags LegendFlags)

@[c: 'ImPlot_SetupMouseText']
fn setup_mouse_text(location Location, flags MouseTextFlags)

@[c: 'ImPlot_SetupFinish']
fn setup_finish()

@[c: 'ImPlot_SetNextAxisLimits']
fn set_next_axis_limits(axis ImAxis, v_min f64, v_max f64, cond Cond)

@[c: 'ImPlot_SetNextAxisLinks']
fn set_next_axis_links(axis ImAxis, link_min &f64, link_max &f64)

@[c: 'ImPlot_SetNextAxisToFit']
fn set_next_axis_to_fit(axis ImAxis)

@[c: 'ImPlot_SetNextAxesLimits']
fn set_next_axes_limits(x_min f64, x_max f64, y_min f64, y_max f64, cond Cond)

@[c: 'ImPlot_SetNextAxesToFit']
fn set_next_axes_to_fit()

@[c: 'ImPlot_PlotLine_FloatPtrInt']
fn plot_line_float_ptr_int(label_id &i8, values &f32, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_doublePtrInt']
fn plot_line_double_ptr_int(label_id &i8, values &f64, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S8PtrInt']
fn plot_line_s8_ptr_int(label_id &i8, values &ImS8, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U8PtrInt']
fn plot_line_u8_ptr_int(label_id &i8, values &ImU8, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S16PtrInt']
fn plot_line_s16_ptr_int(label_id &i8, values &ImS16, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U16PtrInt']
fn plot_line_u16_ptr_int(label_id &i8, values &ImU16, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S32PtrInt']
fn plot_line_s32_ptr_int(label_id &i8, values &ImS32, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U32PtrInt']
fn plot_line_u32_ptr_int(label_id &i8, values &ImU32, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S64PtrInt']
fn plot_line_s64_ptr_int(label_id &i8, values &ImS64, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U64PtrInt']
fn plot_line_u64_ptr_int(label_id &i8, values &ImU64, count int, xscale f64, xstart f64, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_FloatPtrFloatPtr']
fn plot_line_float_ptr_float_ptr(label_id &i8, xs &f32, ys &f32, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_doublePtrdoublePtr']
fn plot_line_double_ptrdouble_ptr(label_id &i8, xs &f64, ys &f64, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S8PtrS8Ptr']
fn plot_line_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U8PtrU8Ptr']
fn plot_line_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S16PtrS16Ptr']
fn plot_line_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U16PtrU16Ptr']
fn plot_line_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S32PtrS32Ptr']
fn plot_line_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U32PtrU32Ptr']
fn plot_line_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_S64PtrS64Ptr']
fn plot_line_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLine_U64PtrU64Ptr']
fn plot_line_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, flags LineFlags, offset int, stride int)

@[c: 'ImPlot_PlotLineG']
fn plot_line_g(label_id &i8, getter Point_getter, data voidptr, count int, flags LineFlags)

// custom generation
@[c: 'ImPlot_PlotScatter_FloatPtrInt']
fn plot_scatter_float_ptr_int(label_id &i8, values &f32, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_doublePtrInt']
fn plot_scatter_double_ptr_int(label_id &i8, values &f64, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S8PtrInt']
fn plot_scatter_s8_ptr_int(label_id &i8, values &ImS8, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U8PtrInt']
fn plot_scatter_u8_ptr_int(label_id &i8, values &ImU8, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S16PtrInt']
fn plot_scatter_s16_ptr_int(label_id &i8, values &ImS16, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U16PtrInt']
fn plot_scatter_u16_ptr_int(label_id &i8, values &ImU16, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S32PtrInt']
fn plot_scatter_s32_ptr_int(label_id &i8, values &ImS32, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U32PtrInt']
fn plot_scatter_u32_ptr_int(label_id &i8, values &ImU32, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S64PtrInt']
fn plot_scatter_s64_ptr_int(label_id &i8, values &ImS64, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U64PtrInt']
fn plot_scatter_u64_ptr_int(label_id &i8, values &ImU64, count int, xscale f64, xstart f64, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_FloatPtrFloatPtr']
fn plot_scatter_float_ptr_float_ptr(label_id &i8, xs &f32, ys &f32, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_doublePtrdoublePtr']
fn plot_scatter_double_ptrdouble_ptr(label_id &i8, xs &f64, ys &f64, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S8PtrS8Ptr']
fn plot_scatter_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U8PtrU8Ptr']
fn plot_scatter_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S16PtrS16Ptr']
fn plot_scatter_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U16PtrU16Ptr']
fn plot_scatter_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S32PtrS32Ptr']
fn plot_scatter_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U32PtrU32Ptr']
fn plot_scatter_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_S64PtrS64Ptr']
fn plot_scatter_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatter_U64PtrU64Ptr']
fn plot_scatter_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, flags ScatterFlags, offset int, stride int)

@[c: 'ImPlot_PlotScatterG']
fn plot_scatter_g(label_id &i8, getter Point_getter, data voidptr, count int, flags ScatterFlags)

// custom generation
@[c: 'ImPlot_PlotStairs_FloatPtrInt']
fn plot_stairs_float_ptr_int(label_id &i8, values &f32, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_doublePtrInt']
fn plot_stairs_double_ptr_int(label_id &i8, values &f64, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S8PtrInt']
fn plot_stairs_s8_ptr_int(label_id &i8, values &ImS8, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U8PtrInt']
fn plot_stairs_u8_ptr_int(label_id &i8, values &ImU8, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S16PtrInt']
fn plot_stairs_s16_ptr_int(label_id &i8, values &ImS16, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U16PtrInt']
fn plot_stairs_u16_ptr_int(label_id &i8, values &ImU16, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S32PtrInt']
fn plot_stairs_s32_ptr_int(label_id &i8, values &ImS32, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U32PtrInt']
fn plot_stairs_u32_ptr_int(label_id &i8, values &ImU32, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S64PtrInt']
fn plot_stairs_s64_ptr_int(label_id &i8, values &ImS64, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U64PtrInt']
fn plot_stairs_u64_ptr_int(label_id &i8, values &ImU64, count int, xscale f64, xstart f64, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_FloatPtrFloatPtr']
fn plot_stairs_float_ptr_float_ptr(label_id &i8, xs &f32, ys &f32, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_doublePtrdoublePtr']
fn plot_stairs_double_ptrdouble_ptr(label_id &i8, xs &f64, ys &f64, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S8PtrS8Ptr']
fn plot_stairs_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U8PtrU8Ptr']
fn plot_stairs_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S16PtrS16Ptr']
fn plot_stairs_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U16PtrU16Ptr']
fn plot_stairs_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S32PtrS32Ptr']
fn plot_stairs_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U32PtrU32Ptr']
fn plot_stairs_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_S64PtrS64Ptr']
fn plot_stairs_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairs_U64PtrU64Ptr']
fn plot_stairs_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, flags StairsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStairsG']
fn plot_stairs_g(label_id &i8, getter Point_getter, data voidptr, count int, flags StairsFlags)

// custom generation
@[c: 'ImPlot_PlotShaded_FloatPtrInt']
fn plot_shaded_float_ptr_int(label_id &i8, values &f32, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_doublePtrInt']
fn plot_shaded_double_ptr_int(label_id &i8, values &f64, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S8PtrInt']
fn plot_shaded_s8_ptr_int(label_id &i8, values &ImS8, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U8PtrInt']
fn plot_shaded_u8_ptr_int(label_id &i8, values &ImU8, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S16PtrInt']
fn plot_shaded_s16_ptr_int(label_id &i8, values &ImS16, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U16PtrInt']
fn plot_shaded_u16_ptr_int(label_id &i8, values &ImU16, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S32PtrInt']
fn plot_shaded_s32_ptr_int(label_id &i8, values &ImS32, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U32PtrInt']
fn plot_shaded_u32_ptr_int(label_id &i8, values &ImU32, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S64PtrInt']
fn plot_shaded_s64_ptr_int(label_id &i8, values &ImS64, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U64PtrInt']
fn plot_shaded_u64_ptr_int(label_id &i8, values &ImU64, count int, yref f64, xscale f64, xstart f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_FloatPtrFloatPtrInt']
fn plot_shaded_float_ptr_float_ptr_int(label_id &i8, xs &f32, ys &f32, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_doublePtrdoublePtrInt']
fn plot_shaded_double_ptrdouble_ptr_int(label_id &i8, xs &f64, ys &f64, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S8PtrS8PtrInt']
fn plot_shaded_s8_ptr_s8_ptr_int(label_id &i8, xs &ImS8, ys &ImS8, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U8PtrU8PtrInt']
fn plot_shaded_u8_ptr_u8_ptr_int(label_id &i8, xs &ImU8, ys &ImU8, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S16PtrS16PtrInt']
fn plot_shaded_s16_ptr_s16_ptr_int(label_id &i8, xs &ImS16, ys &ImS16, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U16PtrU16PtrInt']
fn plot_shaded_u16_ptr_u16_ptr_int(label_id &i8, xs &ImU16, ys &ImU16, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S32PtrS32PtrInt']
fn plot_shaded_s32_ptr_s32_ptr_int(label_id &i8, xs &ImS32, ys &ImS32, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U32PtrU32PtrInt']
fn plot_shaded_u32_ptr_u32_ptr_int(label_id &i8, xs &ImU32, ys &ImU32, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S64PtrS64PtrInt']
fn plot_shaded_s64_ptr_s64_ptr_int(label_id &i8, xs &ImS64, ys &ImS64, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U64PtrU64PtrInt']
fn plot_shaded_u64_ptr_u64_ptr_int(label_id &i8, xs &ImU64, ys &ImU64, count int, yref f64, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_FloatPtrFloatPtrFloatPtr']
fn plot_shaded_float_ptr_float_ptr_float_ptr(label_id &i8, xs &f32, ys1 &f32, ys2 &f32, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_doublePtrdoublePtrdoublePtr']
fn plot_shaded_double_ptrdouble_ptrdouble_ptr(label_id &i8, xs &f64, ys1 &f64, ys2 &f64, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S8PtrS8PtrS8Ptr']
fn plot_shaded_s8_ptr_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys1 &ImS8, ys2 &ImS8, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U8PtrU8PtrU8Ptr']
fn plot_shaded_u8_ptr_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys1 &ImU8, ys2 &ImU8, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S16PtrS16PtrS16Ptr']
fn plot_shaded_s16_ptr_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys1 &ImS16, ys2 &ImS16, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U16PtrU16PtrU16Ptr']
fn plot_shaded_u16_ptr_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys1 &ImU16, ys2 &ImU16, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S32PtrS32PtrS32Ptr']
fn plot_shaded_s32_ptr_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys1 &ImS32, ys2 &ImS32, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U32PtrU32PtrU32Ptr']
fn plot_shaded_u32_ptr_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys1 &ImU32, ys2 &ImU32, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_S64PtrS64PtrS64Ptr']
fn plot_shaded_s64_ptr_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys1 &ImS64, ys2 &ImS64, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShaded_U64PtrU64PtrU64Ptr']
fn plot_shaded_u64_ptr_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys1 &ImU64, ys2 &ImU64, count int, flags ShadedFlags, offset int, stride int)

@[c: 'ImPlot_PlotShadedG']
fn plot_shaded_g(label_id &i8, getter1 Point_getter, data1 voidptr, getter2 Point_getter, data2 voidptr, count int, flags ShadedFlags)

// custom generation
@[c: 'ImPlot_PlotBars_FloatPtrInt']
fn plot_bars_float_ptr_int(label_id &i8, values &f32, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_doublePtrInt']
fn plot_bars_double_ptr_int(label_id &i8, values &f64, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S8PtrInt']
fn plot_bars_s8_ptr_int(label_id &i8, values &ImS8, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U8PtrInt']
fn plot_bars_u8_ptr_int(label_id &i8, values &ImU8, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S16PtrInt']
fn plot_bars_s16_ptr_int(label_id &i8, values &ImS16, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U16PtrInt']
fn plot_bars_u16_ptr_int(label_id &i8, values &ImU16, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S32PtrInt']
fn plot_bars_s32_ptr_int(label_id &i8, values &ImS32, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U32PtrInt']
fn plot_bars_u32_ptr_int(label_id &i8, values &ImU32, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S64PtrInt']
fn plot_bars_s64_ptr_int(label_id &i8, values &ImS64, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U64PtrInt']
fn plot_bars_u64_ptr_int(label_id &i8, values &ImU64, count int, bar_size f64, shift f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_FloatPtrFloatPtr']
fn plot_bars_float_ptr_float_ptr(label_id &i8, xs &f32, ys &f32, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_doublePtrdoublePtr']
fn plot_bars_double_ptrdouble_ptr(label_id &i8, xs &f64, ys &f64, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S8PtrS8Ptr']
fn plot_bars_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U8PtrU8Ptr']
fn plot_bars_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S16PtrS16Ptr']
fn plot_bars_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U16PtrU16Ptr']
fn plot_bars_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S32PtrS32Ptr']
fn plot_bars_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U32PtrU32Ptr']
fn plot_bars_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_S64PtrS64Ptr']
fn plot_bars_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBars_U64PtrU64Ptr']
fn plot_bars_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, bar_size f64, flags BarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotBarsG']
fn plot_bars_g(label_id &i8, getter Point_getter, data voidptr, count int, bar_size f64, flags BarsFlags)

// custom generation
@[c: 'ImPlot_PlotBarGroups_FloatPtr']
fn plot_bar_groups_float_ptr(label_ids &&u8, values &f32, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_doublePtr']
fn plot_bar_groups_double_ptr(label_ids &&u8, values &f64, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_S8Ptr']
fn plot_bar_groups_s8_ptr(label_ids &&u8, values &ImS8, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_U8Ptr']
fn plot_bar_groups_u8_ptr(label_ids &&u8, values &ImU8, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_S16Ptr']
fn plot_bar_groups_s16_ptr(label_ids &&u8, values &ImS16, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_U16Ptr']
fn plot_bar_groups_u16_ptr(label_ids &&u8, values &ImU16, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_S32Ptr']
fn plot_bar_groups_s32_ptr(label_ids &&u8, values &ImS32, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_U32Ptr']
fn plot_bar_groups_u32_ptr(label_ids &&u8, values &ImU32, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_S64Ptr']
fn plot_bar_groups_s64_ptr(label_ids &&u8, values &ImS64, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotBarGroups_U64Ptr']
fn plot_bar_groups_u64_ptr(label_ids &&u8, values &ImU64, item_count int, group_count int, group_size f64, shift f64, flags BarGroupsFlags)

@[c: 'ImPlot_PlotErrorBars_FloatPtrFloatPtrFloatPtrInt']
fn plot_error_bars_float_ptr_float_ptr_float_ptr_int(label_id &i8, xs &f32, ys &f32, err &f32, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_doublePtrdoublePtrdoublePtrInt']
fn plot_error_bars_double_ptrdouble_ptrdouble_ptr_int(label_id &i8, xs &f64, ys &f64, err &f64, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S8PtrS8PtrS8PtrInt']
fn plot_error_bars_s8_ptr_s8_ptr_s8_ptr_int(label_id &i8, xs &ImS8, ys &ImS8, err &ImS8, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U8PtrU8PtrU8PtrInt']
fn plot_error_bars_u8_ptr_u8_ptr_u8_ptr_int(label_id &i8, xs &ImU8, ys &ImU8, err &ImU8, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S16PtrS16PtrS16PtrInt']
fn plot_error_bars_s16_ptr_s16_ptr_s16_ptr_int(label_id &i8, xs &ImS16, ys &ImS16, err &ImS16, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U16PtrU16PtrU16PtrInt']
fn plot_error_bars_u16_ptr_u16_ptr_u16_ptr_int(label_id &i8, xs &ImU16, ys &ImU16, err &ImU16, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S32PtrS32PtrS32PtrInt']
fn plot_error_bars_s32_ptr_s32_ptr_s32_ptr_int(label_id &i8, xs &ImS32, ys &ImS32, err &ImS32, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U32PtrU32PtrU32PtrInt']
fn plot_error_bars_u32_ptr_u32_ptr_u32_ptr_int(label_id &i8, xs &ImU32, ys &ImU32, err &ImU32, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S64PtrS64PtrS64PtrInt']
fn plot_error_bars_s64_ptr_s64_ptr_s64_ptr_int(label_id &i8, xs &ImS64, ys &ImS64, err &ImS64, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U64PtrU64PtrU64PtrInt']
fn plot_error_bars_u64_ptr_u64_ptr_u64_ptr_int(label_id &i8, xs &ImU64, ys &ImU64, err &ImU64, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_FloatPtrFloatPtrFloatPtrFloatPtr']
fn plot_error_bars_float_ptr_float_ptr_float_ptr_float_ptr(label_id &i8, xs &f32, ys &f32, neg &f32, pos &f32, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_doublePtrdoublePtrdoublePtrdoublePtr']
fn plot_error_bars_double_ptrdouble_ptrdouble_ptrdouble_ptr(label_id &i8, xs &f64, ys &f64, neg &f64, pos &f64, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S8PtrS8PtrS8PtrS8Ptr']
fn plot_error_bars_s8_ptr_s8_ptr_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, neg &ImS8, pos &ImS8, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U8PtrU8PtrU8PtrU8Ptr']
fn plot_error_bars_u8_ptr_u8_ptr_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, neg &ImU8, pos &ImU8, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S16PtrS16PtrS16PtrS16Ptr']
fn plot_error_bars_s16_ptr_s16_ptr_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, neg &ImS16, pos &ImS16, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U16PtrU16PtrU16PtrU16Ptr']
fn plot_error_bars_u16_ptr_u16_ptr_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, neg &ImU16, pos &ImU16, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S32PtrS32PtrS32PtrS32Ptr']
fn plot_error_bars_s32_ptr_s32_ptr_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, neg &ImS32, pos &ImS32, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U32PtrU32PtrU32PtrU32Ptr']
fn plot_error_bars_u32_ptr_u32_ptr_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, neg &ImU32, pos &ImU32, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_S64PtrS64PtrS64PtrS64Ptr']
fn plot_error_bars_s64_ptr_s64_ptr_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, neg &ImS64, pos &ImS64, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotErrorBars_U64PtrU64PtrU64PtrU64Ptr']
fn plot_error_bars_u64_ptr_u64_ptr_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, neg &ImU64, pos &ImU64, count int, flags ErrorBarsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_FloatPtrInt']
fn plot_stems_float_ptr_int(label_id &i8, values &f32, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_doublePtrInt']
fn plot_stems_double_ptr_int(label_id &i8, values &f64, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S8PtrInt']
fn plot_stems_s8_ptr_int(label_id &i8, values &ImS8, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U8PtrInt']
fn plot_stems_u8_ptr_int(label_id &i8, values &ImU8, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S16PtrInt']
fn plot_stems_s16_ptr_int(label_id &i8, values &ImS16, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U16PtrInt']
fn plot_stems_u16_ptr_int(label_id &i8, values &ImU16, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S32PtrInt']
fn plot_stems_s32_ptr_int(label_id &i8, values &ImS32, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U32PtrInt']
fn plot_stems_u32_ptr_int(label_id &i8, values &ImU32, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S64PtrInt']
fn plot_stems_s64_ptr_int(label_id &i8, values &ImS64, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U64PtrInt']
fn plot_stems_u64_ptr_int(label_id &i8, values &ImU64, count int, ref f64, scale f64, start f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_FloatPtrFloatPtr']
fn plot_stems_float_ptr_float_ptr(label_id &i8, xs &f32, ys &f32, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_doublePtrdoublePtr']
fn plot_stems_double_ptrdouble_ptr(label_id &i8, xs &f64, ys &f64, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S8PtrS8Ptr']
fn plot_stems_s8_ptr_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U8PtrU8Ptr']
fn plot_stems_u8_ptr_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S16PtrS16Ptr']
fn plot_stems_s16_ptr_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U16PtrU16Ptr']
fn plot_stems_u16_ptr_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S32PtrS32Ptr']
fn plot_stems_s32_ptr_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U32PtrU32Ptr']
fn plot_stems_u32_ptr_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_S64PtrS64Ptr']
fn plot_stems_s64_ptr_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotStems_U64PtrU64Ptr']
fn plot_stems_u64_ptr_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, ref f64, flags StemsFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_FloatPtr']
fn plot_inf_lines_float_ptr(label_id &i8, values &f32, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_doublePtr']
fn plot_inf_lines_double_ptr(label_id &i8, values &f64, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_S8Ptr']
fn plot_inf_lines_s8_ptr(label_id &i8, values &ImS8, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_U8Ptr']
fn plot_inf_lines_u8_ptr(label_id &i8, values &ImU8, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_S16Ptr']
fn plot_inf_lines_s16_ptr(label_id &i8, values &ImS16, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_U16Ptr']
fn plot_inf_lines_u16_ptr(label_id &i8, values &ImU16, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_S32Ptr']
fn plot_inf_lines_s32_ptr(label_id &i8, values &ImS32, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_U32Ptr']
fn plot_inf_lines_u32_ptr(label_id &i8, values &ImU32, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_S64Ptr']
fn plot_inf_lines_s64_ptr(label_id &i8, values &ImS64, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotInfLines_U64Ptr']
fn plot_inf_lines_u64_ptr(label_id &i8, values &ImU64, count int, flags InfLinesFlags, offset int, stride int)

@[c: 'ImPlot_PlotPieChart_FloatPtrPlotFormatter']
fn plot_pie_chart_float_ptr_plot_formatter(label_ids &&u8, values &f32, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_doublePtrPlotFormatter']
fn plot_pie_chart_double_ptr_plot_formatter(label_ids &&u8, values &f64, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S8PtrPlotFormatter']
fn plot_pie_chart_s8_ptr_plot_formatter(label_ids &&u8, values &ImS8, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U8PtrPlotFormatter']
fn plot_pie_chart_u8_ptr_plot_formatter(label_ids &&u8, values &ImU8, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S16PtrPlotFormatter']
fn plot_pie_chart_s16_ptr_plot_formatter(label_ids &&u8, values &ImS16, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U16PtrPlotFormatter']
fn plot_pie_chart_u16_ptr_plot_formatter(label_ids &&u8, values &ImU16, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S32PtrPlotFormatter']
fn plot_pie_chart_s32_ptr_plot_formatter(label_ids &&u8, values &ImS32, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U32PtrPlotFormatter']
fn plot_pie_chart_u32_ptr_plot_formatter(label_ids &&u8, values &ImU32, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S64PtrPlotFormatter']
fn plot_pie_chart_s64_ptr_plot_formatter(label_ids &&u8, values &ImS64, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U64PtrPlotFormatter']
fn plot_pie_chart_u64_ptr_plot_formatter(label_ids &&u8, values &ImU64, count int, x f64, y f64, radius f64, fmt Formatter, fmt_data voidptr, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_FloatPtrStr']
fn plot_pie_chart_float_ptr_str(label_ids &&u8, values &f32, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_doublePtrStr']
fn plot_pie_chart_double_ptr_str(label_ids &&u8, values &f64, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S8PtrStr']
fn plot_pie_chart_s8_ptr_str(label_ids &&u8, values &ImS8, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U8PtrStr']
fn plot_pie_chart_u8_ptr_str(label_ids &&u8, values &ImU8, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S16PtrStr']
fn plot_pie_chart_s16_ptr_str(label_ids &&u8, values &ImS16, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U16PtrStr']
fn plot_pie_chart_u16_ptr_str(label_ids &&u8, values &ImU16, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S32PtrStr']
fn plot_pie_chart_s32_ptr_str(label_ids &&u8, values &ImS32, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U32PtrStr']
fn plot_pie_chart_u32_ptr_str(label_ids &&u8, values &ImU32, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_S64PtrStr']
fn plot_pie_chart_s64_ptr_str(label_ids &&u8, values &ImS64, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotPieChart_U64PtrStr']
fn plot_pie_chart_u64_ptr_str(label_ids &&u8, values &ImU64, count int, x f64, y f64, radius f64, label_fmt &i8, angle0 f64, flags PieChartFlags)

@[c: 'ImPlot_PlotHeatmap_FloatPtr']
fn plot_heatmap_float_ptr(label_id &i8, values &f32, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_doublePtr']
fn plot_heatmap_double_ptr(label_id &i8, values &f64, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_S8Ptr']
fn plot_heatmap_s8_ptr(label_id &i8, values &ImS8, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_U8Ptr']
fn plot_heatmap_u8_ptr(label_id &i8, values &ImU8, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_S16Ptr']
fn plot_heatmap_s16_ptr(label_id &i8, values &ImS16, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_U16Ptr']
fn plot_heatmap_u16_ptr(label_id &i8, values &ImU16, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_S32Ptr']
fn plot_heatmap_s32_ptr(label_id &i8, values &ImS32, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_U32Ptr']
fn plot_heatmap_u32_ptr(label_id &i8, values &ImU32, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_S64Ptr']
fn plot_heatmap_s64_ptr(label_id &i8, values &ImS64, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHeatmap_U64Ptr']
fn plot_heatmap_u64_ptr(label_id &i8, values &ImU64, rows int, cols int, scale_min f64, scale_max f64, label_fmt &i8, bounds_min Point, bounds_max Point, flags HeatmapFlags)

@[c: 'ImPlot_PlotHistogram_FloatPtr']
fn plot_histogram_float_ptr(label_id &i8, values &f32, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_doublePtr']
fn plot_histogram_double_ptr(label_id &i8, values &f64, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_S8Ptr']
fn plot_histogram_s8_ptr(label_id &i8, values &ImS8, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_U8Ptr']
fn plot_histogram_u8_ptr(label_id &i8, values &ImU8, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_S16Ptr']
fn plot_histogram_s16_ptr(label_id &i8, values &ImS16, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_U16Ptr']
fn plot_histogram_u16_ptr(label_id &i8, values &ImU16, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_S32Ptr']
fn plot_histogram_s32_ptr(label_id &i8, values &ImS32, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_U32Ptr']
fn plot_histogram_u32_ptr(label_id &i8, values &ImU32, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_S64Ptr']
fn plot_histogram_s64_ptr(label_id &i8, values &ImS64, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram_U64Ptr']
fn plot_histogram_u64_ptr(label_id &i8, values &ImU64, count int, bins int, bar_scale f64, range Range, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_FloatPtr']
fn plot_histogram2_d_float_ptr(label_id &i8, xs &f32, ys &f32, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_doublePtr']
fn plot_histogram2_d_double_ptr(label_id &i8, xs &f64, ys &f64, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_S8Ptr']
fn plot_histogram2_d_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_U8Ptr']
fn plot_histogram2_d_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_S16Ptr']
fn plot_histogram2_d_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_U16Ptr']
fn plot_histogram2_d_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_S32Ptr']
fn plot_histogram2_d_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_U32Ptr']
fn plot_histogram2_d_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_S64Ptr']
fn plot_histogram2_d_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotHistogram2D_U64Ptr']
fn plot_histogram2_d_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, x_bins int, y_bins int, range Rect, flags HistogramFlags) f64

@[c: 'ImPlot_PlotDigital_FloatPtr']
fn plot_digital_float_ptr(label_id &i8, xs &f32, ys &f32, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_doublePtr']
fn plot_digital_double_ptr(label_id &i8, xs &f64, ys &f64, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_S8Ptr']
fn plot_digital_s8_ptr(label_id &i8, xs &ImS8, ys &ImS8, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_U8Ptr']
fn plot_digital_u8_ptr(label_id &i8, xs &ImU8, ys &ImU8, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_S16Ptr']
fn plot_digital_s16_ptr(label_id &i8, xs &ImS16, ys &ImS16, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_U16Ptr']
fn plot_digital_u16_ptr(label_id &i8, xs &ImU16, ys &ImU16, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_S32Ptr']
fn plot_digital_s32_ptr(label_id &i8, xs &ImS32, ys &ImS32, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_U32Ptr']
fn plot_digital_u32_ptr(label_id &i8, xs &ImU32, ys &ImU32, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_S64Ptr']
fn plot_digital_s64_ptr(label_id &i8, xs &ImS64, ys &ImS64, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigital_U64Ptr']
fn plot_digital_u64_ptr(label_id &i8, xs &ImU64, ys &ImU64, count int, flags DigitalFlags, offset int, stride int)

@[c: 'ImPlot_PlotDigitalG']
fn plot_digital_g(label_id &i8, getter Point_getter, data voidptr, count int, flags DigitalFlags)

// custom generation
@[c: 'ImPlot_PlotImage']
fn plot_image(label_id &i8, user_texture_id ImTextureID, bounds_min Point, bounds_max Point, uv0 ImVec2, uv1 ImVec2, tint_col C.ImVec4, flags ImageFlags)

@[c: 'ImPlot_PlotText']
fn plot_text(text &i8, x f64, y f64, pix_offset ImVec2, flags TextFlags)

@[c: 'ImPlot_PlotDummy']
fn plot_dummy(label_id &i8, flags DummyFlags)

@[c: 'ImPlot_DragPoint']
fn drag_point(id int, x &f64, y &f64, col C.ImVec4, size f32, flags DragToolFlags, out_clicked &bool, out_hovered &bool, held &bool) bool

@[c: 'ImPlot_DragLineX']
fn drag_line_x(id int, x &f64, col C.ImVec4, thickness f32, flags DragToolFlags, out_clicked &bool, out_hovered &bool, held &bool) bool

@[c: 'ImPlot_DragLineY']
fn drag_line_y(id int, y &f64, col C.ImVec4, thickness f32, flags DragToolFlags, out_clicked &bool, out_hovered &bool, held &bool) bool

@[c: 'ImPlot_DragRect']
fn drag_rect(id int, x1 &f64, y1 &f64, x2 &f64, y2 &f64, col C.ImVec4, flags DragToolFlags, out_clicked &bool, out_hovered &bool, held &bool) bool

@[c: 'ImPlot_Annotation_Bool']
fn annotation_bool(x f64, y f64, col C.ImVec4, pix_offset ImVec2, clamp bool, round bool)

@[c: 'ImPlot_Annotation_Str']
@[c2v_variadic]
fn annotation_str(x f64, y f64, col C.ImVec4, pix_offset ImVec2, clamp bool, fmt ...&i8)

@[c: 'ImPlot_AnnotationV']
fn annotation_v(x f64, y f64, col C.ImVec4, pix_offset ImVec2, clamp bool, fmt &i8, args C.va_list)

@[c: 'ImPlot_TagX_Bool']
fn tag_x_bool(x f64, col C.ImVec4, round bool)

@[c: 'ImPlot_TagX_Str']
@[c2v_variadic]
fn tag_x_str(x f64, col C.ImVec4, fmt ...&i8)

@[c: 'ImPlot_TagXV']
fn tag_xv(x f64, col C.ImVec4, fmt &i8, args C.va_list)

@[c: 'ImPlot_TagY_Bool']
fn tag_y_bool(y f64, col C.ImVec4, round bool)

@[c: 'ImPlot_TagY_Str']
@[c2v_variadic]
fn tag_y_str(y f64, col C.ImVec4, fmt ...&i8)

@[c: 'ImPlot_TagYV']
fn tag_yv(y f64, col C.ImVec4, fmt &i8, args C.va_list)

@[c: 'ImPlot_SetAxis']
fn set_axis(axis ImAxis)

@[c: 'ImPlot_SetAxes']
fn set_axes(x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_PixelsToPlot_Vec2']
fn pixels_to_plot_vec2(p_out &Point, pix ImVec2, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_PixelsToPlot_Float']
fn pixels_to_plot_float(p_out &Point, x f32, y f32, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_PlotToPixels_PlotPoInt']
fn plot_to_pixels_plot_po_int(p_out &ImVec2, plt Point, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_PlotToPixels_double']
fn plot_to_pixels_double(p_out &ImVec2, x f64, y f64, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_GetPlotPos']
fn get_plot_pos(p_out &ImVec2)

@[c: 'ImPlot_GetPlotSize']
fn get_plot_size(p_out &ImVec2)

@[c: 'ImPlot_GetPlotMousePos']
fn get_plot_mouse_pos(p_out &Point, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_GetPlotLimits']
fn get_plot_limits(p_out &Rect, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_IsPlotHovered']
fn is_plot_hovered() bool

@[c: 'ImPlot_IsAxisHovered']
fn is_axis_hovered(axis ImAxis) bool

@[c: 'ImPlot_IsSubplotsHovered']
fn is_subplots_hovered() bool

@[c: 'ImPlot_IsPlotSelected']
fn is_plot_selected() bool

@[c: 'ImPlot_GetPlotSelection']
fn get_plot_selection(p_out &Rect, x_axis ImAxis, y_axis ImAxis)

@[c: 'ImPlot_CancelPlotSelection']
fn cancel_plot_selection()

@[c: 'ImPlot_HideNextItem']
fn hide_next_item(hidden bool, cond Cond)

@[c: 'ImPlot_BeginAlignedPlots']
fn begin_aligned_plots(group_id &i8, vertical bool) bool

@[c: 'ImPlot_EndAlignedPlots']
fn end_aligned_plots()

@[c: 'ImPlot_BeginLegendPopup']
fn begin_legend_popup(label_id &i8, mouse_button ImGuiMouseButton) bool

@[c: 'ImPlot_EndLegendPopup']
fn end_legend_popup()

@[c: 'ImPlot_IsLegendEntryHovered']
fn is_legend_entry_hovered(label_id &i8) bool

@[c: 'ImPlot_BeginDragDropTargetPlot']
fn begin_drag_drop_target_plot() bool

@[c: 'ImPlot_BeginDragDropTargetAxis']
fn begin_drag_drop_target_axis(axis ImAxis) bool

@[c: 'ImPlot_BeginDragDropTargetLegend']
fn begin_drag_drop_target_legend() bool

@[c: 'ImPlot_EndDragDropTarget']
fn end_drag_drop_target()

@[c: 'ImPlot_BeginDragDropSourcePlot']
fn begin_drag_drop_source_plot(flags ImGuiDragDropFlags) bool

@[c: 'ImPlot_BeginDragDropSourceAxis']
fn begin_drag_drop_source_axis(axis ImAxis, flags ImGuiDragDropFlags) bool

@[c: 'ImPlot_BeginDragDropSourceItem']
fn begin_drag_drop_source_item(label_id &i8, flags ImGuiDragDropFlags) bool

@[c: 'ImPlot_EndDragDropSource']
fn end_drag_drop_source()

@[c: 'ImPlot_GetStyle']
fn get_style() &Style

@[c: 'ImPlot_StyleColorsAuto']
fn style_colors_auto(dst &Style)

@[c: 'ImPlot_StyleColorsClassic']
fn style_colors_classic(dst &Style)

@[c: 'ImPlot_StyleColorsDark']
fn style_colors_dark(dst &Style)

@[c: 'ImPlot_StyleColorsLight']
fn style_colors_light(dst &Style)

@[c: 'ImPlot_PushStyleColor_U32']
fn push_style_color_u32(idx Col, col ImU32)

@[c: 'ImPlot_PushStyleColor_Vec4']
fn push_style_color_vec4(idx Col, col C.ImVec4)

@[c: 'ImPlot_PopStyleColor']
fn pop_style_color(count int)

@[c: 'ImPlot_PushStyleVar_Float']
fn push_style_var_float(idx StyleVar, val f32)

@[c: 'ImPlot_PushStyleVar_Int']
fn push_style_var_int(idx StyleVar, val int)

@[c: 'ImPlot_PushStyleVar_Vec2']
fn push_style_var_vec2(idx StyleVar, val ImVec2)

@[c: 'ImPlot_PopStyleVar']
fn pop_style_var(count int)

@[c: 'ImPlot_SetNextLineStyle']
fn set_next_line_style(col C.ImVec4, weight f32)

@[c: 'ImPlot_SetNextFillStyle']
fn set_next_fill_style(col C.ImVec4, alpha_mod f32)

@[c: 'ImPlot_SetNextMarkerStyle']
fn set_next_marker_style(marker Marker, size f32, fill C.ImVec4, weight f32, outline C.ImVec4)

@[c: 'ImPlot_SetNextErrorBarStyle']
fn set_next_error_bar_style(col C.ImVec4, size f32, weight f32)

@[c: 'ImPlot_GetLastItemColor']
fn get_last_item_color(p_out &C.ImVec4)

@[c: 'ImPlot_GetStyleColorName']
fn get_style_color_name(idx Col) &i8

@[c: 'ImPlot_GetMarkerName']
fn get_marker_name(idx Marker) &i8

@[c: 'ImPlot_AddColormap_Vec4Ptr']
fn add_colormap_vec4_ptr(name &i8, cols &C.ImVec4, size int, qual bool) Colormap

@[c: 'ImPlot_AddColormap_U32Ptr']
fn add_colormap_u32_ptr(name &i8, cols &ImU32, size int, qual bool) Colormap

@[c: 'ImPlot_GetColormapCount']
fn get_colormap_count() int

@[c: 'ImPlot_GetColormapName']
fn get_colormap_name(cmap Colormap) &i8

@[c: 'ImPlot_GetColormapIndex']
fn get_colormap_index(name &i8) Colormap

@[c: 'ImPlot_PushColormap_PlotColormap']
fn push_colormap_plot_colormap(cmap Colormap)

@[c: 'ImPlot_PushColormap_Str']
fn push_colormap_str(name &i8)

@[c: 'ImPlot_PopColormap']
fn pop_colormap(count int)

@[c: 'ImPlot_NextColormapColor']
fn next_colormap_color(p_out &C.ImVec4)

@[c: 'ImPlot_GetColormapSize']
fn get_colormap_size(cmap Colormap) int

@[c: 'ImPlot_GetColormapColor']
fn get_colormap_color(p_out &C.ImVec4, idx int, cmap Colormap)

@[c: 'ImPlot_SampleColormap']
fn sample_colormap(p_out &C.ImVec4, t f32, cmap Colormap)

@[c: 'ImPlot_ColormapScale']
fn colormap_scale(label &i8, scale_min f64, scale_max f64, size ImVec2, format &i8, flags ColormapScaleFlags, cmap Colormap)

@[c: 'ImPlot_ColormapSlider']
fn colormap_slider(label &i8, t &f32, out &C.ImVec4, format &i8, cmap Colormap) bool

@[c: 'ImPlot_ColormapButton']
fn colormap_button(label &i8, size ImVec2, cmap Colormap) bool

@[c: 'ImPlot_BustColorCache']
fn bust_color_cache(plot_title_id &i8)

@[c: 'ImPlot_GetInputMap']
fn get_input_map() &InputMap

@[c: 'ImPlot_MapInputDefault']
fn map_input_default(dst &InputMap)

@[c: 'ImPlot_MapInputReverse']
fn map_input_reverse(dst &InputMap)

@[c: 'ImPlot_ItemIcon_Vec4']
fn item_icon_vec4(col C.ImVec4)

@[c: 'ImPlot_ItemIcon_U32']
fn item_icon_u32(col ImU32)

@[c: 'ImPlot_ColormapIcon']
fn colormap_icon(cmap Colormap)

@[c: 'ImPlot_GetPlotDrawList']
fn get_plot_draw_list() &ImDrawList

@[c: 'ImPlot_PushPlotClipRect']
fn push_plot_clip_rect(expand f32)

@[c: 'ImPlot_PopPlotClipRect']
fn pop_plot_clip_rect()

@[c: 'ImPlot_ShowStyleSelector']
fn show_style_selector(label &i8) bool

@[c: 'ImPlot_ShowColormapSelector']
fn show_colormap_selector(label &i8) bool

@[c: 'ImPlot_ShowInputMapSelector']
fn show_input_map_selector(label &i8) bool

@[c: 'ImPlot_ShowStyleEditor']
fn show_style_editor(ref &Style)

@[c: 'ImPlot_ShowUserGuide']
fn show_user_guide()

@[c: 'ImPlot_ShowMetricsWindow']
fn show_metrics_window(p_popen &bool)

@[c: 'ImPlot_ShowDemoWindow']
fn show_demo_window(p_open &bool)

@[c: 'ImPlot_ImLog10_Float']
fn im_log10_float(x f32) f32

@[c: 'ImPlot_ImLog10_double']
fn im_log10_double(x f64) f64

@[c: 'ImPlot_ImSinh_Float']
fn im_sinh_float(x f32) f32

@[c: 'ImPlot_ImSinh_double']
fn im_sinh_double(x f64) f64

@[c: 'ImPlot_ImAsinh_Float']
fn im_asinh_float(x f32) f32

@[c: 'ImPlot_ImAsinh_double']
fn im_asinh_double(x f64) f64

@[c: 'ImPlot_ImRemap_Float']
fn im_remap_float(x f32, x0 f32, x1 f32, y0 f32, y1 f32) f32

@[c: 'ImPlot_ImRemap_double']
fn im_remap_double(x f64, x0 f64, x1 f64, y0 f64, y1 f64) f64

@[c: 'ImPlot_ImRemap_S8']
fn im_remap_s8(x ImS8, x0 ImS8, x1 ImS8, y0 ImS8, y1 ImS8) ImS8

@[c: 'ImPlot_ImRemap_U8']
fn im_remap_u8(x ImU8, x0 ImU8, x1 ImU8, y0 ImU8, y1 ImU8) ImU8

@[c: 'ImPlot_ImRemap_S16']
fn im_remap_s16(x ImS16, x0 ImS16, x1 ImS16, y0 ImS16, y1 ImS16) ImS16

@[c: 'ImPlot_ImRemap_U16']
fn im_remap_u16(x ImU16, x0 ImU16, x1 ImU16, y0 ImU16, y1 ImU16) ImU16

@[c: 'ImPlot_ImRemap_S32']
fn im_remap_s32(x ImS32, x0 ImS32, x1 ImS32, y0 ImS32, y1 ImS32) ImS32

@[c: 'ImPlot_ImRemap_U32']
fn im_remap_u32(x ImU32, x0 ImU32, x1 ImU32, y0 ImU32, y1 ImU32) ImU32

@[c: 'ImPlot_ImRemap_S64']
fn im_remap_s64(x ImS64, x0 ImS64, x1 ImS64, y0 ImS64, y1 ImS64) ImS64

@[c: 'ImPlot_ImRemap_U64']
fn im_remap_u64(x ImU64, x0 ImU64, x1 ImU64, y0 ImU64, y1 ImU64) ImU64

@[c: 'ImPlot_ImRemap01_Float']
fn im_remap01_float(x f32, x0 f32, x1 f32) f32

@[c: 'ImPlot_ImRemap01_double']
fn im_remap01_double(x f64, x0 f64, x1 f64) f64

@[c: 'ImPlot_ImRemap01_S8']
fn im_remap01_s8(x ImS8, x0 ImS8, x1 ImS8) ImS8

@[c: 'ImPlot_ImRemap01_U8']
fn im_remap01_u8(x ImU8, x0 ImU8, x1 ImU8) ImU8

@[c: 'ImPlot_ImRemap01_S16']
fn im_remap01_s16(x ImS16, x0 ImS16, x1 ImS16) ImS16

@[c: 'ImPlot_ImRemap01_U16']
fn im_remap01_u16(x ImU16, x0 ImU16, x1 ImU16) ImU16

@[c: 'ImPlot_ImRemap01_S32']
fn im_remap01_s32(x ImS32, x0 ImS32, x1 ImS32) ImS32

@[c: 'ImPlot_ImRemap01_U32']
fn im_remap01_u32(x ImU32, x0 ImU32, x1 ImU32) ImU32

@[c: 'ImPlot_ImRemap01_S64']
fn im_remap01_s64(x ImS64, x0 ImS64, x1 ImS64) ImS64

@[c: 'ImPlot_ImRemap01_U64']
fn im_remap01_u64(x ImU64, x0 ImU64, x1 ImU64) ImU64

@[c: 'ImPlot_ImPosMod']
fn im_pos_mod(l int, r int) int

@[c: 'ImPlot_ImNan']
fn im_nan(val f64) bool

@[c: 'ImPlot_ImNanOrInf']
fn im_nan_or_inf(val f64) bool

@[c: 'ImPlot_ImConstrainNan']
fn im_constrain_nan(val f64) f64

@[c: 'ImPlot_ImConstrainInf']
fn im_constrain_inf(val f64) f64

@[c: 'ImPlot_ImConstrainLog']
fn im_constrain_log(val f64) f64

@[c: 'ImPlot_ImConstrainTime']
fn im_constrain_time(val f64) f64

@[c: 'ImPlot_ImAlmostEqual']
fn im_almost_equal(v1 f64, v2 f64, ulp int) bool

@[c: 'ImPlot_ImMinArray_FloatPtr']
fn im_min_array_float_ptr(values &f32, count int) f32

@[c: 'ImPlot_ImMinArray_doublePtr']
fn im_min_array_double_ptr(values &f64, count int) f64

@[c: 'ImPlot_ImMinArray_S8Ptr']
fn im_min_array_s8_ptr(values &ImS8, count int) ImS8

@[c: 'ImPlot_ImMinArray_U8Ptr']
fn im_min_array_u8_ptr(values &ImU8, count int) ImU8

@[c: 'ImPlot_ImMinArray_S16Ptr']
fn im_min_array_s16_ptr(values &ImS16, count int) ImS16

@[c: 'ImPlot_ImMinArray_U16Ptr']
fn im_min_array_u16_ptr(values &ImU16, count int) ImU16

@[c: 'ImPlot_ImMinArray_S32Ptr']
fn im_min_array_s32_ptr(values &ImS32, count int) ImS32

@[c: 'ImPlot_ImMinArray_U32Ptr']
fn im_min_array_u32_ptr(values &ImU32, count int) ImU32

@[c: 'ImPlot_ImMinArray_S64Ptr']
fn im_min_array_s64_ptr(values &ImS64, count int) ImS64

@[c: 'ImPlot_ImMinArray_U64Ptr']
fn im_min_array_u64_ptr(values &ImU64, count int) ImU64

@[c: 'ImPlot_ImMaxArray_FloatPtr']
fn im_max_array_float_ptr(values &f32, count int) f32

@[c: 'ImPlot_ImMaxArray_doublePtr']
fn im_max_array_double_ptr(values &f64, count int) f64

@[c: 'ImPlot_ImMaxArray_S8Ptr']
fn im_max_array_s8_ptr(values &ImS8, count int) ImS8

@[c: 'ImPlot_ImMaxArray_U8Ptr']
fn im_max_array_u8_ptr(values &ImU8, count int) ImU8

@[c: 'ImPlot_ImMaxArray_S16Ptr']
fn im_max_array_s16_ptr(values &ImS16, count int) ImS16

@[c: 'ImPlot_ImMaxArray_U16Ptr']
fn im_max_array_u16_ptr(values &ImU16, count int) ImU16

@[c: 'ImPlot_ImMaxArray_S32Ptr']
fn im_max_array_s32_ptr(values &ImS32, count int) ImS32

@[c: 'ImPlot_ImMaxArray_U32Ptr']
fn im_max_array_u32_ptr(values &ImU32, count int) ImU32

@[c: 'ImPlot_ImMaxArray_S64Ptr']
fn im_max_array_s64_ptr(values &ImS64, count int) ImS64

@[c: 'ImPlot_ImMaxArray_U64Ptr']
fn im_max_array_u64_ptr(values &ImU64, count int) ImU64

@[c: 'ImPlot_ImMinMaxArray_FloatPtr']
fn im_min_max_array_float_ptr(values &f32, count int, min_out &f32, max_out &f32)

@[c: 'ImPlot_ImMinMaxArray_doublePtr']
fn im_min_max_array_double_ptr(values &f64, count int, min_out &f64, max_out &f64)

@[c: 'ImPlot_ImMinMaxArray_S8Ptr']
fn im_min_max_array_s8_ptr(values &ImS8, count int, min_out &ImS8, max_out &ImS8)

@[c: 'ImPlot_ImMinMaxArray_U8Ptr']
fn im_min_max_array_u8_ptr(values &ImU8, count int, min_out &ImU8, max_out &ImU8)

@[c: 'ImPlot_ImMinMaxArray_S16Ptr']
fn im_min_max_array_s16_ptr(values &ImS16, count int, min_out &ImS16, max_out &ImS16)

@[c: 'ImPlot_ImMinMaxArray_U16Ptr']
fn im_min_max_array_u16_ptr(values &ImU16, count int, min_out &ImU16, max_out &ImU16)

@[c: 'ImPlot_ImMinMaxArray_S32Ptr']
fn im_min_max_array_s32_ptr(values &ImS32, count int, min_out &ImS32, max_out &ImS32)

@[c: 'ImPlot_ImMinMaxArray_U32Ptr']
fn im_min_max_array_u32_ptr(values &ImU32, count int, min_out &ImU32, max_out &ImU32)

@[c: 'ImPlot_ImMinMaxArray_S64Ptr']
fn im_min_max_array_s64_ptr(values &ImS64, count int, min_out &ImS64, max_out &ImS64)

@[c: 'ImPlot_ImMinMaxArray_U64Ptr']
fn im_min_max_array_u64_ptr(values &ImU64, count int, min_out &ImU64, max_out &ImU64)

@[c: 'ImPlot_ImSum_FloatPtr']
fn im_sum_float_ptr(values &f32, count int) f32

@[c: 'ImPlot_ImSum_doublePtr']
fn im_sum_double_ptr(values &f64, count int) f64

@[c: 'ImPlot_ImSum_S8Ptr']
fn im_sum_s8_ptr(values &ImS8, count int) ImS8

@[c: 'ImPlot_ImSum_U8Ptr']
fn im_sum_u8_ptr(values &ImU8, count int) ImU8

@[c: 'ImPlot_ImSum_S16Ptr']
fn im_sum_s16_ptr(values &ImS16, count int) ImS16

@[c: 'ImPlot_ImSum_U16Ptr']
fn im_sum_u16_ptr(values &ImU16, count int) ImU16

@[c: 'ImPlot_ImSum_S32Ptr']
fn im_sum_s32_ptr(values &ImS32, count int) ImS32

@[c: 'ImPlot_ImSum_U32Ptr']
fn im_sum_u32_ptr(values &ImU32, count int) ImU32

@[c: 'ImPlot_ImSum_S64Ptr']
fn im_sum_s64_ptr(values &ImS64, count int) ImS64

@[c: 'ImPlot_ImSum_U64Ptr']
fn im_sum_u64_ptr(values &ImU64, count int) ImU64

@[c: 'ImPlot_ImMean_FloatPtr']
fn im_mean_float_ptr(values &f32, count int) f64

@[c: 'ImPlot_ImMean_doublePtr']
fn im_mean_double_ptr(values &f64, count int) f64

@[c: 'ImPlot_ImMean_S8Ptr']
fn im_mean_s8_ptr(values &ImS8, count int) f64

@[c: 'ImPlot_ImMean_U8Ptr']
fn im_mean_u8_ptr(values &ImU8, count int) f64

@[c: 'ImPlot_ImMean_S16Ptr']
fn im_mean_s16_ptr(values &ImS16, count int) f64

@[c: 'ImPlot_ImMean_U16Ptr']
fn im_mean_u16_ptr(values &ImU16, count int) f64

@[c: 'ImPlot_ImMean_S32Ptr']
fn im_mean_s32_ptr(values &ImS32, count int) f64

@[c: 'ImPlot_ImMean_U32Ptr']
fn im_mean_u32_ptr(values &ImU32, count int) f64

@[c: 'ImPlot_ImMean_S64Ptr']
fn im_mean_s64_ptr(values &ImS64, count int) f64

@[c: 'ImPlot_ImMean_U64Ptr']
fn im_mean_u64_ptr(values &ImU64, count int) f64

@[c: 'ImPlot_ImStdDev_FloatPtr']
fn im_std_dev_float_ptr(values &f32, count int) f64

@[c: 'ImPlot_ImStdDev_doublePtr']
fn im_std_dev_double_ptr(values &f64, count int) f64

@[c: 'ImPlot_ImStdDev_S8Ptr']
fn im_std_dev_s8_ptr(values &ImS8, count int) f64

@[c: 'ImPlot_ImStdDev_U8Ptr']
fn im_std_dev_u8_ptr(values &ImU8, count int) f64

@[c: 'ImPlot_ImStdDev_S16Ptr']
fn im_std_dev_s16_ptr(values &ImS16, count int) f64

@[c: 'ImPlot_ImStdDev_U16Ptr']
fn im_std_dev_u16_ptr(values &ImU16, count int) f64

@[c: 'ImPlot_ImStdDev_S32Ptr']
fn im_std_dev_s32_ptr(values &ImS32, count int) f64

@[c: 'ImPlot_ImStdDev_U32Ptr']
fn im_std_dev_u32_ptr(values &ImU32, count int) f64

@[c: 'ImPlot_ImStdDev_S64Ptr']
fn im_std_dev_s64_ptr(values &ImS64, count int) f64

@[c: 'ImPlot_ImStdDev_U64Ptr']
fn im_std_dev_u64_ptr(values &ImU64, count int) f64

@[c: 'ImPlot_ImMixU32']
fn im_mix_u32(a ImU32, b ImU32, s ImU32) ImU32

@[c: 'ImPlot_ImLerpU32']
fn im_lerp_u32(colors &ImU32, size int, t f32) ImU32

@[c: 'ImPlot_ImAlphaU32']
fn im_alpha_u32(col ImU32, alpha f32) ImU32

@[c: 'ImPlot_ImOverlaps_Float']
fn im_overlaps_float(min_a f32, max_a f32, min_b f32, max_b f32) bool

@[c: 'ImPlot_ImOverlaps_double']
fn im_overlaps_double(min_a f64, max_a f64, min_b f64, max_b f64) bool

@[c: 'ImPlot_ImOverlaps_S8']
fn im_overlaps_s8(min_a ImS8, max_a ImS8, min_b ImS8, max_b ImS8) bool

@[c: 'ImPlot_ImOverlaps_U8']
fn im_overlaps_u8(min_a ImU8, max_a ImU8, min_b ImU8, max_b ImU8) bool

@[c: 'ImPlot_ImOverlaps_S16']
fn im_overlaps_s16(min_a ImS16, max_a ImS16, min_b ImS16, max_b ImS16) bool

@[c: 'ImPlot_ImOverlaps_U16']
fn im_overlaps_u16(min_a ImU16, max_a ImU16, min_b ImU16, max_b ImU16) bool

@[c: 'ImPlot_ImOverlaps_S32']
fn im_overlaps_s32(min_a ImS32, max_a ImS32, min_b ImS32, max_b ImS32) bool

@[c: 'ImPlot_ImOverlaps_U32']
fn im_overlaps_u32(min_a ImU32, max_a ImU32, min_b ImU32, max_b ImU32) bool

@[c: 'ImPlot_ImOverlaps_S64']
fn im_overlaps_s64(min_a ImS64, max_a ImS64, min_b ImS64, max_b ImS64) bool

@[c: 'ImPlot_ImOverlaps_U64']
fn im_overlaps_u64(min_a ImU64, max_a ImU64, min_b ImU64, max_b ImU64) bool

@[c: 'ImPlotDateTimeSpec_ImPlotDateTimeSpec_Nil']
fn date_time_spec_im_plot_date_time_spec_nil() &DateTimeSpec

@[c: 'ImPlotDateTimeSpec_destroy']
fn date_time_spec_destroy(self &DateTimeSpec)

@[c: 'ImPlotDateTimeSpec_ImPlotDateTimeSpec_PlotDateFmt']
fn date_time_spec_im_plot_date_time_spec_plot_date_fmt(date_fmt DateFmt, time_fmt TimeFmt, use_24_hr_clk bool, use_iso_8601 bool) &DateTimeSpec

@[c: 'ImPlotTime_ImPlotTime_Nil']
fn time_im_plot_time_nil() &Time

@[c: 'ImPlotTime_destroy']
fn time_destroy(self &Time)

@[c: 'ImPlotTime_ImPlotTime_time_t']
fn time_im_plot_time_time_t(s C.time_t, us int) &Time

@[c: 'ImPlotTime_RollOver']
fn time_roll_over(self &Time)

@[c: 'ImPlotTime_ToDouble']
fn time_to_double(self &Time) f64

@[c: 'ImPlotTime_FromDouble']
fn time_from_double(p_out &Time, t f64)

@[c: 'ImPlotColormapData_ImPlotColormapData']
fn colormap_data_im_plot_colormap_data() &ColormapData

@[c: 'ImPlotColormapData_destroy']
fn colormap_data_destroy(self &ColormapData)

@[c: 'ImPlotColormapData_Append']
fn colormap_data_append(self &ColormapData, name &i8, keys &ImU32, count int, qual bool) int

@[c: 'ImPlotColormapData__AppendTable']
fn colormap_data__append_table(self &ColormapData, cmap Colormap)

@[c: 'ImPlotColormapData_RebuildTables']
fn colormap_data_rebuild_tables(self &ColormapData)

@[c: 'ImPlotColormapData_IsQual']
fn colormap_data_is_qual(self &ColormapData, cmap Colormap) bool

@[c: 'ImPlotColormapData_GetName']
fn colormap_data_get_name(self &ColormapData, cmap Colormap) &i8

@[c: 'ImPlotColormapData_GetIndex']
fn colormap_data_get_index(self &ColormapData, name &i8) Colormap

@[c: 'ImPlotColormapData_GetKeys']
fn colormap_data_get_keys(self &ColormapData, cmap Colormap) &ImU32

@[c: 'ImPlotColormapData_GetKeyCount']
fn colormap_data_get_key_count(self &ColormapData, cmap Colormap) int

@[c: 'ImPlotColormapData_GetKeyColor']
fn colormap_data_get_key_color(self &ColormapData, cmap Colormap, idx int) ImU32

@[c: 'ImPlotColormapData_SetKeyColor']
fn colormap_data_set_key_color(self &ColormapData, cmap Colormap, idx int, value ImU32)

@[c: 'ImPlotColormapData_GetTable']
fn colormap_data_get_table(self &ColormapData, cmap Colormap) &ImU32

@[c: 'ImPlotColormapData_GetTableSize']
fn colormap_data_get_table_size(self &ColormapData, cmap Colormap) int

@[c: 'ImPlotColormapData_GetTableColor']
fn colormap_data_get_table_color(self &ColormapData, cmap Colormap, idx int) ImU32

@[c: 'ImPlotColormapData_LerpTable']
fn colormap_data_lerp_table(self &ColormapData, cmap Colormap, t f32) ImU32

@[c: 'ImPlotPointError_ImPlotPointError']
fn point_error_im_plot_point_error(x f64, y f64, neg f64, pos f64) &PointError

@[c: 'ImPlotPointError_destroy']
fn point_error_destroy(self &PointError)

@[c: 'ImPlotAnnotation_ImPlotAnnotation']
fn annotation_im_plot_annotation() &Annotation

@[c: 'ImPlotAnnotation_destroy']
fn annotation_destroy(self &Annotation)

@[c: 'ImPlotAnnotationCollection_ImPlotAnnotationCollection']
fn annotation_collection_im_plot_annotation_collection() &AnnotationCollection

@[c: 'ImPlotAnnotationCollection_destroy']
fn annotation_collection_destroy(self &AnnotationCollection)

@[c: 'ImPlotAnnotationCollection_AppendV']
fn annotation_collection_append_v(self &AnnotationCollection, pos ImVec2, off ImVec2, bg ImU32, fg ImU32, clamp bool, fmt &i8, args C.va_list)

@[c: 'ImPlotAnnotationCollection_Append']
@[c2v_variadic]
fn annotation_collection_append(self &AnnotationCollection, pos ImVec2, off ImVec2, bg ImU32, fg ImU32, clamp bool, fmt ...&i8)

@[c: 'ImPlotAnnotationCollection_GetText']
fn annotation_collection_get_text(self &AnnotationCollection, idx int) &i8

@[c: 'ImPlotAnnotationCollection_Reset']
fn annotation_collection_reset(self &AnnotationCollection)

@[c: 'ImPlotTagCollection_ImPlotTagCollection']
fn tag_collection_im_plot_tag_collection() &TagCollection

@[c: 'ImPlotTagCollection_destroy']
fn tag_collection_destroy(self &TagCollection)

@[c: 'ImPlotTagCollection_AppendV']
fn tag_collection_append_v(self &TagCollection, axis ImAxis, value f64, bg ImU32, fg ImU32, fmt &i8, args C.va_list)

@[c: 'ImPlotTagCollection_Append']
@[c2v_variadic]
fn tag_collection_append(self &TagCollection, axis ImAxis, value f64, bg ImU32, fg ImU32, fmt ...&i8)

@[c: 'ImPlotTagCollection_GetText']
fn tag_collection_get_text(self &TagCollection, idx int) &i8

@[c: 'ImPlotTagCollection_Reset']
fn tag_collection_reset(self &TagCollection)

@[c: 'ImPlotTick_ImPlotTick']
fn tick_im_plot_tick(value f64, major bool, level int, show_label bool) &Tick

@[c: 'ImPlotTick_destroy']
fn tick_destroy(self &Tick)

@[c: 'ImPlotTicker_ImPlotTicker']
fn ticker_im_plot_ticker() &Ticker

@[c: 'ImPlotTicker_destroy']
fn ticker_destroy(self &Ticker)

@[c: 'ImPlotTicker_AddTick_doubleStr']
fn ticker_add_tick_double_str(self &Ticker, value f64, major bool, level int, show_label bool, label &i8) &Tick

@[c: 'ImPlotTicker_AddTick_doublePlotFormatter']
fn ticker_add_tick_double_plot_formatter(self &Ticker, value f64, major bool, level int, show_label bool, formatter Formatter, data voidptr) &Tick

@[c: 'ImPlotTicker_AddTick_PlotTick']
fn ticker_add_tick_plot_tick(self &Ticker, tick Tick) &Tick

@[c: 'ImPlotTicker_GetText_Int']
fn ticker_get_text_int(self &Ticker, idx int) &i8

@[c: 'ImPlotTicker_GetText_PlotTick']
fn ticker_get_text_plot_tick(self &Ticker, tick Tick) &i8

@[c: 'ImPlotTicker_OverrideSizeLate']
fn ticker_override_size_late(self &Ticker, size ImVec2)

@[c: 'ImPlotTicker_Reset']
fn ticker_reset(self &Ticker)

@[c: 'ImPlotTicker_TickCount']
fn ticker_tick_count(self &Ticker) int

@[c: 'ImPlotAxis_ImPlotAxis']
fn axis_im_plot_axis() &Axis

@[c: 'ImPlotAxis_destroy']
fn axis_destroy(self &Axis)

@[c: 'ImPlotAxis_Reset']
fn axis_reset(self &Axis)

@[c: 'ImPlotAxis_SetMin']
fn axis_set_min(self &Axis, _min f64, force bool) bool

@[c: 'ImPlotAxis_SetMax']
fn axis_set_max(self &Axis, _max f64, force bool) bool

@[c: 'ImPlotAxis_SetRange_double']
fn axis_set_range_double(self &Axis, v1 f64, v2 f64)

@[c: 'ImPlotAxis_SetRange_PlotRange']
fn axis_set_range_plot_range(self &Axis, range Range)

@[c: 'ImPlotAxis_SetAspect']
fn axis_set_aspect(self &Axis, unit_per_pix f64)

@[c: 'ImPlotAxis_PixelSize']
fn axis_pixel_size(self &Axis) f32

@[c: 'ImPlotAxis_GetAspect']
fn axis_get_aspect(self &Axis) f64

@[c: 'ImPlotAxis_Constrain']
fn axis_constrain(self &Axis)

@[c: 'ImPlotAxis_UpdateTransformCache']
fn axis_update_transform_cache(self &Axis)

@[c: 'ImPlotAxis_PlotToPixels']
fn axis_plot_to_pixels(self &Axis, plt f64) f32

@[c: 'ImPlotAxis_PixelsToPlot']
fn axis_pixels_to_plot(self &Axis, pix f32) f64

@[c: 'ImPlotAxis_ExtendFit']
fn axis_extend_fit(self &Axis, v f64)

@[c: 'ImPlotAxis_ExtendFitWith']
fn axis_extend_fit_with(self &Axis, alt &Axis, v f64, v_alt f64)

@[c: 'ImPlotAxis_ApplyFit']
fn axis_apply_fit(self &Axis, padding f32)

@[c: 'ImPlotAxis_HasLabel']
fn axis_has_label(self &Axis) bool

@[c: 'ImPlotAxis_HasGridLines']
fn axis_has_grid_lines(self &Axis) bool

@[c: 'ImPlotAxis_HasTickLabels']
fn axis_has_tick_labels(self &Axis) bool

@[c: 'ImPlotAxis_HasTickMarks']
fn axis_has_tick_marks(self &Axis) bool

@[c: 'ImPlotAxis_WillRender']
fn axis_will_render(self &Axis) bool

@[c: 'ImPlotAxis_IsOpposite']
fn axis_is_opposite(self &Axis) bool

@[c: 'ImPlotAxis_IsInverted']
fn axis_is_inverted(self &Axis) bool

@[c: 'ImPlotAxis_IsForeground']
fn axis_is_foreground(self &Axis) bool

@[c: 'ImPlotAxis_IsAutoFitting']
fn axis_is_auto_fitting(self &Axis) bool

@[c: 'ImPlotAxis_CanInitFit']
fn axis_can_init_fit(self &Axis) bool

@[c: 'ImPlotAxis_IsRangeLocked']
fn axis_is_range_locked(self &Axis) bool

@[c: 'ImPlotAxis_IsLockedMin']
fn axis_is_locked_min(self &Axis) bool

@[c: 'ImPlotAxis_IsLockedMax']
fn axis_is_locked_max(self &Axis) bool

@[c: 'ImPlotAxis_IsLocked']
fn axis_is_locked(self &Axis) bool

@[c: 'ImPlotAxis_IsInputLockedMin']
fn axis_is_input_locked_min(self &Axis) bool

@[c: 'ImPlotAxis_IsInputLockedMax']
fn axis_is_input_locked_max(self &Axis) bool

@[c: 'ImPlotAxis_IsInputLocked']
fn axis_is_input_locked(self &Axis) bool

@[c: 'ImPlotAxis_HasMenus']
fn axis_has_menus(self &Axis) bool

@[c: 'ImPlotAxis_IsPanLocked']
fn axis_is_pan_locked(self &Axis, increasing bool) bool

@[c: 'ImPlotAxis_PushLinks']
fn axis_push_links(self &Axis)

@[c: 'ImPlotAxis_PullLinks']
fn axis_pull_links(self &Axis)

@[c: 'ImPlotAlignmentData_ImPlotAlignmentData']
fn alignment_data_im_plot_alignment_data() &AlignmentData

@[c: 'ImPlotAlignmentData_destroy']
fn alignment_data_destroy(self &AlignmentData)

@[c: 'ImPlotAlignmentData_Begin']
fn alignment_data_begin(self &AlignmentData)

@[c: 'ImPlotAlignmentData_Update']
fn alignment_data_update(self &AlignmentData, pad_a &f32, pad_b &f32, delta_a &f32, delta_b &f32)

@[c: 'ImPlotAlignmentData_End']
fn alignment_data_end(self &AlignmentData)

@[c: 'ImPlotAlignmentData_Reset']
fn alignment_data_reset(self &AlignmentData)

@[c: 'ImPlotItem_ImPlotItem']
fn item_im_plot_item() &Item

@[c: 'ImPlotItem_destroy']
fn item_destroy(self &Item)

@[c: 'ImPlotLegend_ImPlotLegend']
fn legend_im_plot_legend() &Legend

@[c: 'ImPlotLegend_destroy']
fn legend_destroy(self &Legend)

@[c: 'ImPlotLegend_Reset']
fn legend_reset(self &Legend)

@[c: 'ImPlotItemGroup_ImPlotItemGroup']
fn item_group_im_plot_item_group() &ItemGroup

@[c: 'ImPlotItemGroup_destroy']
fn item_group_destroy(self &ItemGroup)

@[c: 'ImPlotItemGroup_GetItemCount']
fn item_group_get_item_count(self &ItemGroup) int

@[c: 'ImPlotItemGroup_GetItemID']
fn item_group_get_item_id(self &ItemGroup, label_id &i8) ImGuiID

@[c: 'ImPlotItemGroup_GetItem_ID']
fn item_group_get_item_id_vdup0(self &ItemGroup, id ImGuiID) &Item

@[c: 'ImPlotItemGroup_GetItem_Str']
fn item_group_get_item_str(self &ItemGroup, label_id &i8) &Item

@[c: 'ImPlotItemGroup_GetOrAddItem']
fn item_group_get_or_add_item(self &ItemGroup, id ImGuiID) &Item

@[c: 'ImPlotItemGroup_GetItemByIndex']
fn item_group_get_item_by_index(self &ItemGroup, i int) &Item

@[c: 'ImPlotItemGroup_GetItemIndex']
fn item_group_get_item_index(self &ItemGroup, item &Item) int

@[c: 'ImPlotItemGroup_GetLegendCount']
fn item_group_get_legend_count(self &ItemGroup) int

@[c: 'ImPlotItemGroup_GetLegendItem']
fn item_group_get_legend_item(self &ItemGroup, i int) &Item

@[c: 'ImPlotItemGroup_GetLegendLabel']
fn item_group_get_legend_label(self &ItemGroup, i int) &i8

@[c: 'ImPlotItemGroup_Reset']
fn item_group_reset(self &ItemGroup)

@[c: 'ImPlotPlot_ImPlotPlot']
fn plot_im_plot_plot() &Plot

@[c: 'ImPlotPlot_destroy']
fn plot_destroy(self &Plot)

@[c: 'ImPlotPlot_IsInputLocked']
fn plot_is_input_locked(self &Plot) bool

@[c: 'ImPlotPlot_ClearTextBuffer']
fn plot_clear_text_buffer(self &Plot)

@[c: 'ImPlotPlot_SetTitle']
fn plot_set_title(self &Plot, title &i8)

@[c: 'ImPlotPlot_HasTitle']
fn plot_has_title(self &Plot) bool

@[c: 'ImPlotPlot_GetTitle']
fn plot_get_title(self &Plot) &i8

@[c: 'ImPlotPlot_XAxis_Nil']
fn plot_xa_xis_nil(self &Plot, i int) &Axis

@[c: 'ImPlotPlot_XAxis__const']
fn plot_xa_xis__const(self &Plot, i int) &Axis

@[c: 'ImPlotPlot_YAxis_Nil']
fn plot_ya_xis_nil(self &Plot, i int) &Axis

@[c: 'ImPlotPlot_YAxis__const']
fn plot_ya_xis__const(self &Plot, i int) &Axis

@[c: 'ImPlotPlot_EnabledAxesX']
fn plot_enabled_axes_x(self &Plot) int

@[c: 'ImPlotPlot_EnabledAxesY']
fn plot_enabled_axes_y(self &Plot) int

@[c: 'ImPlotPlot_SetAxisLabel']
fn plot_set_axis_label(self &Plot, axis &Axis, label &i8)

@[c: 'ImPlotPlot_GetAxisLabel']
fn plot_get_axis_label(self &Plot, axis Axis) &i8

@[c: 'ImPlotSubplot_ImPlotSubplot']
fn subplot_im_plot_subplot() &Subplot

@[c: 'ImPlotSubplot_destroy']
fn subplot_destroy(self &Subplot)

@[c: 'ImPlotNextPlotData_ImPlotNextPlotData']
fn next_plot_data_im_plot_next_plot_data() &NextPlotData

@[c: 'ImPlotNextPlotData_destroy']
fn next_plot_data_destroy(self &NextPlotData)

@[c: 'ImPlotNextPlotData_Reset']
fn next_plot_data_reset(self &NextPlotData)

@[c: 'ImPlotNextItemData_ImPlotNextItemData']
fn next_item_data_im_plot_next_item_data() &NextItemData

@[c: 'ImPlotNextItemData_destroy']
fn next_item_data_destroy(self &NextItemData)

@[c: 'ImPlotNextItemData_Reset']
fn next_item_data_reset(self &NextItemData)

@[c: 'ImPlot_Initialize']
fn initialize(ctx &Context)

@[c: 'ImPlot_ResetCtxForNextPlot']
fn reset_ctx_for_next_plot(ctx &Context)

@[c: 'ImPlot_ResetCtxForNextAlignedPlots']
fn reset_ctx_for_next_aligned_plots(ctx &Context)

@[c: 'ImPlot_ResetCtxForNextSubplot']
fn reset_ctx_for_next_subplot(ctx &Context)

@[c: 'ImPlot_GetPlot']
fn get_plot(title &i8) &Plot

@[c: 'ImPlot_GetCurrentPlot']
fn get_current_plot() &Plot

@[c: 'ImPlot_BustPlotCache']
fn bust_plot_cache()

@[c: 'ImPlot_ShowPlotContextMenu']
fn show_plot_context_menu(plot &Plot)

@[c: 'ImPlot_SetupLock']
fn setup_lock()

@[c: 'ImPlot_SubplotNextCell']
fn subplot_next_cell()

@[c: 'ImPlot_ShowSubplotsContextMenu']
fn show_subplots_context_menu(subplot &Subplot)

@[c: 'ImPlot_BeginItem']
fn begin_item(label_id &i8, flags ItemFlags, recolor_from Col) bool

@[c: 'ImPlot_EndItem']
fn end_item()

@[c: 'ImPlot_RegisterOrGetItem']
fn register_or_get_item(label_id &i8, flags ItemFlags, just_created &bool) &Item

@[c: 'ImPlot_GetItem']
fn get_item(label_id &i8) &Item

@[c: 'ImPlot_GetCurrentItem']
fn get_current_item() &Item

@[c: 'ImPlot_BustItemCache']
fn bust_item_cache()

@[c: 'ImPlot_AnyAxesInputLocked']
fn any_axes_input_locked(axes &Axis, count int) bool

@[c: 'ImPlot_AllAxesInputLocked']
fn all_axes_input_locked(axes &Axis, count int) bool

@[c: 'ImPlot_AnyAxesHeld']
fn any_axes_held(axes &Axis, count int) bool

@[c: 'ImPlot_AnyAxesHovered']
fn any_axes_hovered(axes &Axis, count int) bool

@[c: 'ImPlot_FitThisFrame']
fn fit_this_frame() bool

@[c: 'ImPlot_FitPointX']
fn fit_point_x(x f64)

@[c: 'ImPlot_FitPointY']
fn fit_point_y(y f64)

@[c: 'ImPlot_FitPoint']
fn fit_point(p Point)

@[c: 'ImPlot_RangesOverlap']
fn ranges_overlap(r1 Range, r2 Range) bool

@[c: 'ImPlot_ShowAxisContextMenu']
fn show_axis_context_menu(axis &Axis, equal_axis &Axis, time_allowed bool)

@[c: 'ImPlot_GetLocationPos']
fn get_location_pos(p_out &ImVec2, outer_rect C.ImRect, inner_size ImVec2, location Location, pad ImVec2)

@[c: 'ImPlot_CalcLegendSize']
fn calc_legend_size(p_out &ImVec2, items &ItemGroup, pad ImVec2, spacing ImVec2, vertical bool)

@[c: 'ImPlot_ClampLegendRect']
fn clamp_legend_rect(legend_rect &C.ImRect, outer_rect C.ImRect, pad ImVec2) bool

@[c: 'ImPlot_ShowLegendEntries']
fn show_legend_entries(items &ItemGroup, legend_bb C.ImRect, interactable bool, pad ImVec2, spacing ImVec2, vertical bool, draw_list &ImDrawList) bool

@[c: 'ImPlot_ShowAltLegend']
fn show_alt_legend(title_id &i8, vertical bool, size ImVec2, interactable bool)

@[c: 'ImPlot_ShowLegendContextMenu']
fn show_legend_context_menu(legend &Legend, visible bool) bool

@[c: 'ImPlot_LabelAxisValue']
fn label_axis_value(axis Axis, value f64, buff &i8, size int, round bool)

@[c: 'ImPlot_GetItemData']
fn get_item_data() &NextItemData

@[c: 'ImPlot_IsColorAuto_Vec4']
fn is_color_auto_vec4(col C.ImVec4) bool

@[c: 'ImPlot_IsColorAuto_PlotCol']
fn is_color_auto_plot_col(idx Col) bool

@[c: 'ImPlot_GetAutoColor']
fn get_auto_color(p_out &C.ImVec4, idx Col)

@[c: 'ImPlot_GetStyleColorVec4']
fn get_style_color_vec4(p_out &C.ImVec4, idx Col)

@[c: 'ImPlot_GetStyleColorU32']
fn get_style_color_u32(idx Col) ImU32

@[c: 'ImPlot_AddTextVertical']
fn add_text_vertical(draw_list &ImDrawList, pos ImVec2, col ImU32, text_begin &i8, text_end &i8)

@[c: 'ImPlot_AddTextCentered']
fn add_text_centered(draw_list &ImDrawList, top_center ImVec2, col ImU32, text_begin &i8, text_end &i8)

@[c: 'ImPlot_CalcTextSizeVertical']
fn calc_text_size_vertical(p_out &ImVec2, text &i8)

@[c: 'ImPlot_CalcTextColor_Vec4']
fn calc_text_color_vec4(bg C.ImVec4) ImU32

@[c: 'ImPlot_CalcTextColor_U32']
fn calc_text_color_u32(bg ImU32) ImU32

@[c: 'ImPlot_CalcHoverColor']
fn calc_hover_color(col ImU32) ImU32

@[c: 'ImPlot_ClampLabelPos']
fn clamp_label_pos(p_out &ImVec2, pos ImVec2, size ImVec2, min ImVec2, max ImVec2)

@[c: 'ImPlot_GetColormapColorU32']
fn get_colormap_color_u32(idx int, cmap Colormap) ImU32

@[c: 'ImPlot_NextColormapColorU32']
fn next_colormap_color_u32() ImU32

@[c: 'ImPlot_SampleColormapU32']
fn sample_colormap_u32(t f32, cmap Colormap) ImU32

@[c: 'ImPlot_RenderColorBar']
fn render_color_bar(colors &ImU32, size int, draw_list &ImDrawList, bounds C.ImRect, vert bool, reversed bool, continuous bool)

@[c: 'ImPlot_NiceNum']
fn nice_num(x f64, round bool) f64

@[c: 'ImPlot_OrderOfMagnitude']
fn order_of_magnitude(val f64) int

@[c: 'ImPlot_OrderToPrecision']
fn order_to_precision(order int) int

@[c: 'ImPlot_Precision']
fn precision(val f64) int

@[c: 'ImPlot_RoundTo']
fn round_to(val f64, prec int) f64

@[c: 'ImPlot_Intersection']
fn intersection(p_out &ImVec2, a1 ImVec2, a2 ImVec2, b1 ImVec2, b2 ImVec2)

@[c: 'ImPlot_FillRange_Vector_Float_Ptr']
fn fill_range_vector_float_ptr(buffer &ImVector_float, n int, vmin f32, vmax f32)

@[c: 'ImPlot_FillRange_Vector_double_Ptr']
fn fill_range_vector_double_ptr(buffer &ImVector_double, n int, vmin f64, vmax f64)

@[c: 'ImPlot_FillRange_Vector_S8_Ptr']
fn fill_range_vector_s8_ptr(buffer &ImVector_ImS8, n int, vmin ImS8, vmax ImS8)

@[c: 'ImPlot_FillRange_Vector_U8_Ptr']
fn fill_range_vector_u8_ptr(buffer &ImVector_ImU8, n int, vmin ImU8, vmax ImU8)

@[c: 'ImPlot_FillRange_Vector_S16_Ptr']
fn fill_range_vector_s16_ptr(buffer &ImVector_ImS16, n int, vmin ImS16, vmax ImS16)

@[c: 'ImPlot_FillRange_Vector_U16_Ptr']
fn fill_range_vector_u16_ptr(buffer &ImVector_ImU16, n int, vmin ImU16, vmax ImU16)

@[c: 'ImPlot_FillRange_Vector_S32_Ptr']
fn fill_range_vector_s32_ptr(buffer &ImVector_ImS32, n int, vmin ImS32, vmax ImS32)

@[c: 'ImPlot_FillRange_Vector_U32_Ptr']
fn fill_range_vector_u32_ptr(buffer &ImVector_ImU32, n int, vmin ImU32, vmax ImU32)

@[c: 'ImPlot_FillRange_Vector_S64_Ptr']
fn fill_range_vector_s64_ptr(buffer &ImVector_ImS64, n int, vmin ImS64, vmax ImS64)

@[c: 'ImPlot_FillRange_Vector_U64_Ptr']
fn fill_range_vector_u64_ptr(buffer &ImVector_ImU64, n int, vmin ImU64, vmax ImU64)

@[c: 'ImPlot_CalculateBins_FloatPtr']
fn calculate_bins_float_ptr(values &f32, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_doublePtr']
fn calculate_bins_double_ptr(values &f64, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_S8Ptr']
fn calculate_bins_s8_ptr(values &ImS8, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_U8Ptr']
fn calculate_bins_u8_ptr(values &ImU8, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_S16Ptr']
fn calculate_bins_s16_ptr(values &ImS16, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_U16Ptr']
fn calculate_bins_u16_ptr(values &ImU16, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_S32Ptr']
fn calculate_bins_s32_ptr(values &ImS32, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_U32Ptr']
fn calculate_bins_u32_ptr(values &ImU32, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_S64Ptr']
fn calculate_bins_s64_ptr(values &ImS64, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_CalculateBins_U64Ptr']
fn calculate_bins_u64_ptr(values &ImU64, count int, meth Bin, range Range, bins_out &int, width_out &f64)

@[c: 'ImPlot_IsLeapYear']
fn is_leap_year(year int) bool

@[c: 'ImPlot_GetDaysInMonth']
fn get_days_in_month(year int, month int) int

@[c: 'ImPlot_MkGmtTime']
fn mk_gmt_time(p_out &Time, ptm &C.tm)

@[c: 'ImPlot_GetGmtTime']
fn get_gmt_time(t Time, ptm &C.tm) &C.tm

@[c: 'ImPlot_MkLocTime']
fn mk_loc_time(p_out &Time, ptm &C.tm)

@[c: 'ImPlot_GetLocTime']
fn get_loc_time(t Time, ptm &C.tm) &C.tm

@[c: 'ImPlot_MkTime']
fn mk_time(p_out &Time, ptm &C.tm)

@[c: 'ImPlot_GetTime']
fn get_time(t Time, ptm &C.tm) &C.tm

@[c: 'ImPlot_MakeTime']
fn make_time(p_out &Time, year int, month int, day int, hour int, min int, sec int, us int)

@[c: 'ImPlot_GetYear']
fn get_year(t Time) int

@[c: 'ImPlot_GetMonth']
fn get_month(t Time) int

@[c: 'ImPlot_AddTime']
fn add_time(p_out &Time, t Time, unit TimeUnit, count int)

@[c: 'ImPlot_FloorTime']
fn floor_time(p_out &Time, t Time, unit TimeUnit)

@[c: 'ImPlot_CeilTime']
fn ceil_time(p_out &Time, t Time, unit TimeUnit)

@[c: 'ImPlot_RoundTime']
fn round_time(p_out &Time, t Time, unit TimeUnit)

@[c: 'ImPlot_CombineDateTime']
fn combine_date_time(p_out &Time, date_part Time, time_part Time)

@[c: 'ImPlot_Now']
fn now(p_out &Time)

@[c: 'ImPlot_Today']
fn today(p_out &Time)

@[c: 'ImPlot_FormatTime']
fn format_time(t Time, buffer &i8, size int, fmt TimeFmt, use_24_hr_clk bool) int

@[c: 'ImPlot_FormatDate']
fn format_date(t Time, buffer &i8, size int, fmt DateFmt, use_iso_8601 bool) int

@[c: 'ImPlot_FormatDateTime']
fn format_date_time(t Time, buffer &i8, size int, fmt DateTimeSpec) int

@[c: 'ImPlot_ShowDatePicker']
fn show_date_picker(id &i8, level &int, t &Time, t1 &Time, t2 &Time) bool

@[c: 'ImPlot_ShowTimePicker']
fn show_time_picker(id &i8, t &Time) bool

@[c: 'ImPlot_TransformForward_Log10']
fn transform_forward_log10(v f64, noname1 voidptr) f64

@[c: 'ImPlot_TransformInverse_Log10']
fn transform_inverse_log10(v f64, noname1 voidptr) f64

@[c: 'ImPlot_TransformForward_SymLog']
fn transform_forward_sym_log(v f64, noname1 voidptr) f64

@[c: 'ImPlot_TransformInverse_SymLog']
fn transform_inverse_sym_log(v f64, noname1 voidptr) f64

@[c: 'ImPlot_TransformForward_Logit']
fn transform_forward_logit(v f64, noname1 voidptr) f64

@[c: 'ImPlot_TransformInverse_Logit']
fn transform_inverse_logit(v f64, noname1 voidptr) f64

@[c: 'ImPlot_Formatter_Default']
fn formatter_default(value f64, buff &i8, size int, data voidptr) int

@[c: 'ImPlot_Formatter_Logit']
fn formatter_logit(value f64, buff &i8, size int, noname1 voidptr) int

@[c: 'ImPlot_Formatter_Time']
fn formatter_time(noname1 f64, buff &i8, size int, data voidptr) int

@[c: 'ImPlot_Locator_Default']
fn locator_default(ticker &Ticker, range Range, pixels f32, vertical bool, formatter Formatter, formatter_data voidptr)

@[c: 'ImPlot_Locator_Time']
fn locator_time(ticker &Ticker, range Range, pixels f32, vertical bool, formatter Formatter, formatter_data voidptr)

@[c: 'ImPlot_Locator_Log10']
fn locator_log10(ticker &Ticker, range Range, pixels f32, vertical bool, formatter Formatter, formatter_data voidptr)

@[c: 'ImPlot_Locator_SymLog']
fn locator_sym_log(ticker &Ticker, range Range, pixels f32, vertical bool, formatter Formatter, formatter_data voidptr)

// CIMGUIPLOT_INCLUDED
