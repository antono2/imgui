@[translated]
module imgui

#flag -I @VMODROOT/include
#include <cimgui.h>
#flag -DCIMGUI_DEFINE_ENUMS_AND_STRUCTS
#flag -DIMGUI_USE_WCHAR32

pub const version = '1.91.9b'
pub const version_num = 19191

pub type C.ImGuiDockNodeSettings = voidptr
pub type C.ImGuiTabBar = voidptr
pub type C.ImGuiSizeCallback = voidptr
pub type C.ImGuiSelectionExternalStorage = voidptr
pub type C.ImGuiInputTextCallback = voidptr
pub type C.ImBitVector = voidptr
pub type C.ImGuiIDStackTool = voidptr
pub type C.ImWchar = voidptr
pub type C.ImGuiInputEvent = voidptr
pub type C.ImGuiLocEntry = voidptr
pub type C.ImVec4 = voidptr
pub type C.ImGuiDockRequest = voidptr
pub type C.ImRect = voidptr
pub type C.va_list = voidptr
pub type C.ImGuiTextFilter = voidptr

// This file is automatically generated by int(generator.lua) from https://int(github.com)/cimgui/cimgui
// based on int(imgui.h) file version "1.91.9b" 19191 from Dear ImGui https://int(github.com)/ocornut/imgui
// with int(imgui_internal.h) api
// with int(imgui_freetype.h) api
// docking branch
// typedef unsigned long long ImU64;
struct ImVector_const_charPtr {
	size     int
	capacity int
	data     &&u8
}

type ID = u32
type ImS8 = i8
type ImU8 = u8
type ImS16 = i16
type ImU16 = u16
type ImS32 = int
type ImU32 = u32
type ImS64 = i64
type ImU64 = i64
type Col = int
type Cond = int
type DataType = int
type MouseButton = int
type MouseCursor = int
type StyleVar = int
type TableBgTarget = int
type ImDrawFlags = int
type ImDrawListFlags = int
type ImFontAtlasFlags = int
type BackendFlags = int
type ButtonFlags = int
type ChildFlags = int
type ColorEditFlags = int
type ConfigFlags = int
type ComboFlags = int
type DockNodeFlags = int
type DragDropFlags = int
type FocusedFlags = int
type HoveredFlags = int
type InputFlags = int
type InputTextFlags = int
type ItemFlags = int
type KeyChord = int
type PopupFlags = int
type MultiSelectFlags = int
type SelectableFlags = int
type SliderFlags = int
type ImGuiTabBarFlags = int
type TabItemFlags = int
type TableFlags = int
type TableColumnFlags = int
type TableRowFlags = int
type TreeNodeFlags = int
type ViewportFlags = int
type WindowFlags = int
type ImWchar32 = u32
type ImWchar16 = u16
type SelectionUserData = i64
type MemAllocFunc = fn (usize, voidptr) voidptr

type MemFreeFunc = fn (voidptr, voidptr)

struct ImVec2 {
	x f32
	y f32
}

struct ImTextureID {
	x f32
	y f32
	z f32
	w f32
}

enum WindowFlags_ {
	none                        = 0
	no_title_bar                = 1 << 0
	no_resize                   = 1 << 1
	no_move                     = 1 << 2
	no_scrollbar                = 1 << 3
	no_scroll_with_mouse        = 1 << 4
	no_collapse                 = 1 << 5
	always_auto_resize          = 1 << 6
	no_background               = 1 << 7
	no_saved_settings           = 1 << 8
	no_mouse_inputs             = 1 << 9
	menu_bar                    = 1 << 10
	horizontal_scrollbar        = 1 << 11
	no_focus_on_appearing       = 1 << 12
	no_bring_to_front_on_focus  = 1 << 13
	always_vertical_scrollbar   = 1 << 14
	always_horizontal_scrollbar = 1 << 15
	no_nav_inputs               = 1 << 16
	no_nav_focus                = 1 << 17
	unsaved_document            = 1 << 18
	no_docking                  = 1 << 19
	no_nav                      = 1 << 16 | 1 << 17
	no_decoration               = 1 << 0 | 1 << 1 | 1 << 3 | 1 << 5
	no_inputs                   = 1 << 9 | 1 << 16 | 1 << 17
	dock_node_host              = 1 << 23
	child_window                = 1 << 24
	tooltip                     = 1 << 25
	popup                       = 1 << 26
	modal                       = 1 << 27
	child_menu                  = 1 << 28
}

enum ChildFlags_ {
	none                      = 0
	borders                   = 1 << 0
	always_use_window_padding = 1 << 1
	resize_x                  = 1 << 2
	resize_y                  = 1 << 3
	auto_resize_x             = 1 << 4
	auto_resize_y             = 1 << 5
	always_auto_resize        = 1 << 6
	frame_style               = 1 << 7
	nav_flattened             = 1 << 8
}

enum ItemFlags_ {
	none                 = 0
	no_tab_stop          = 1 << 0
	no_nav               = 1 << 1
	no_nav_default_focus = 1 << 2
	button_repeat        = 1 << 3
	auto_close_popups    = 1 << 4
	allow_duplicate_id   = 1 << 5
}

enum InputTextFlags_ {
	none                    = 0
	chars_decimal           = 1 << 0
	chars_hexadecimal       = 1 << 1
	chars_scientific        = 1 << 2
	chars_uppercase         = 1 << 3
	chars_no_blank          = 1 << 4
	allow_tab_input         = 1 << 5
	enter_returns_true      = 1 << 6
	escape_clears_all       = 1 << 7
	ctrl_enter_for_new_line = 1 << 8
	read_only               = 1 << 9
	password                = 1 << 10
	always_overwrite        = 1 << 11
	auto_select_all         = 1 << 12
	parse_empty_ref_val     = 1 << 13
	display_empty_ref_val   = 1 << 14
	no_horizontal_scroll    = 1 << 15
	no_undo_redo            = 1 << 16
	elide_left              = 1 << 17
	callback_completion     = 1 << 18
	callback_history        = 1 << 19
	callback_always         = 1 << 20
	callback_char_filter    = 1 << 21
	callback_resize         = 1 << 22
	callback_edit           = 1 << 23
}

enum TreeNodeFlags_ {
	none                     = 0
	selected                 = 1 << 0
	framed                   = 1 << 1
	allow_overlap            = 1 << 2
	no_tree_push_on_open     = 1 << 3
	no_auto_open_on_log      = 1 << 4
	default_open             = 1 << 5
	open_on_double_click     = 1 << 6
	open_on_arrow            = 1 << 7
	leaf                     = 1 << 8
	bullet                   = 1 << 9
	frame_padding            = 1 << 10
	span_avail_width         = 1 << 11
	span_full_width          = 1 << 12
	span_label_width         = 1 << 13
	span_all_columns         = 1 << 14
	label_span_all_columns   = 1 << 15
	nav_left_jumps_back_here = 1 << 17
	collapsing_header        = 1 << 1 | 1 << 3 | 1 << 4
}

enum PopupFlags_ {
	none                        = 0
	mouse_button_left           = 0
	mouse_button_right          = 1
	mouse_button_middle         = 2
	mouse_button_mask_          = 31
	mouse_button_default_       = 1
	no_reopen                   = 1 << 5
	no_open_over_existing_popup = 1 << 7
	no_open_over_items          = 1 << 8
	any_popup_id                = 1 << 10
	any_popup_level             = 1 << 11
	any_popup                   = 1 << 10 | 1 << 11
}

enum SelectableFlags_ {
	none                 = 0
	no_auto_close_popups = 1 << 0
	span_all_columns     = 1 << 1
	allow_double_click   = 1 << 2
	disabled             = 1 << 3
	allow_overlap        = 1 << 4
	highlight            = 1 << 5
}

enum ComboFlags_ {
	none              = 0
	popup_align_left  = 1 << 0
	height_small      = 1 << 1
	height_regular    = 1 << 2
	height_large      = 1 << 3
	height_largest    = 1 << 4
	no_arrow_button   = 1 << 5
	no_preview        = 1 << 6
	width_fit_preview = 1 << 7
	height_mask_      = 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4
}

enum ImGuiTabBarFlags_ {
	none                              = 0
	reorderable                       = 1 << 0
	auto_select_new_tabs              = 1 << 1
	tab_list_popup_button             = 1 << 2
	no_close_with_middle_mouse_button = 1 << 3
	no_tab_list_scrolling_buttons     = 1 << 4
	no_tooltip                        = 1 << 5
	draw_selected_overline            = 1 << 6
	fitting_policy_resize_down        = 1 << 7
	fitting_policy_scroll             = 1 << 8
	fitting_policy_mask_              = 1 << 7 | 1 << 8
	fitting_policy_default_           = 1 << 7
}

enum TabItemFlags_ {
	none                              = 0
	unsaved_document                  = 1 << 0
	set_selected                      = 1 << 1
	no_close_with_middle_mouse_button = 1 << 2
	no_push_id                        = 1 << 3
	no_tooltip                        = 1 << 4
	no_reorder                        = 1 << 5
	leading                           = 1 << 6
	trailing                          = 1 << 7
	no_assumed_closure                = 1 << 8
}

enum FocusedFlags_ {
	none                   = 0
	child_windows          = 1 << 0
	root_window            = 1 << 1
	any_window             = 1 << 2
	no_popup_hierarchy     = 1 << 3
	dock_hierarchy         = 1 << 4
	root_and_child_windows = 1 << 1 | 1 << 0
}

enum HoveredFlags_ {
	none                              = 0
	child_windows                     = 1 << 0
	root_window                       = 1 << 1
	any_window                        = 1 << 2
	no_popup_hierarchy                = 1 << 3
	dock_hierarchy                    = 1 << 4
	allow_when_blocked_by_popup       = 1 << 5
	allow_when_blocked_by_active_item = 1 << 7
	allow_when_overlapped_by_item     = 1 << 8
	allow_when_overlapped_by_window   = 1 << 9
	allow_when_disabled               = 1 << 10
	no_nav_override                   = 1 << 11
	allow_when_overlapped             = 1 << 8 | 1 << 9
	rect_only                         = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9
	root_and_child_windows            = 1 << 1 | 1 << 0
	for_tooltip                       = 1 << 12
	stationary                        = 1 << 13
	delay_none                        = 1 << 14
	delay_short                       = 1 << 15
	delay_normal                      = 1 << 16
	no_shared_delay                   = 1 << 17
}

enum DockNodeFlags_ {
	none                         = 0
	keep_alive_only              = 1 << 0
	no_docking_over_central_node = 1 << 2
	passthru_central_node        = 1 << 3
	no_docking_split             = 1 << 4
	no_resize                    = 1 << 5
	auto_hide_tab_bar            = 1 << 6
	no_undocking                 = 1 << 7
}

enum DragDropFlags_ {
	none                          = 0
	source_no_preview_tooltip     = 1 << 0
	source_no_disable_hover       = 1 << 1
	source_no_hold_to_open_others = 1 << 2
	source_allow_null_id          = 1 << 3
	source_extern                 = 1 << 4
	payload_auto_expire           = 1 << 5
	payload_no_cross_context      = 1 << 6
	payload_no_cross_process      = 1 << 7
	accept_before_delivery        = 1 << 10
	accept_no_draw_default_rect   = 1 << 11
	accept_no_preview_tooltip     = 1 << 12
	accept_peek_only              = 1 << 10 | 1 << 11
}

enum DataType_ {
	s8
	u8
	s16
	u16
	s32
	u32
	s64
	u64
	float
	double
	bool
	string
	count
}

enum Dir {
	none  = -1
	left  = 0
	right = 1
	up    = 2
	down  = 3
	count = 4
}

enum SortDirection {
	none       = 0
	ascending  = 1
	descending = 2
}

enum Key {
	none                   = 0
	named_begin            = 512
	tab                    = 512
	left_arrow             = 513
	right_arrow            = 514
	up_arrow               = 515
	down_arrow             = 516
	page_up                = 517
	page_down              = 518
	home                   = 519
	end                    = 520
	insert                 = 521
	delete                 = 522
	backspace              = 523
	space                  = 524
	enter                  = 525
	escape                 = 526
	left_ctrl              = 527
	left_shift             = 528
	left_alt               = 529
	left_super             = 530
	right_ctrl             = 531
	right_shift            = 532
	right_alt              = 533
	right_super            = 534
	menu                   = 535
	_0                     = 536
	_1                     = 537
	_2                     = 538
	_3                     = 539
	_4                     = 540
	_5                     = 541
	_6                     = 542
	_7                     = 543
	_8                     = 544
	_9                     = 545
	a                      = 546
	b                      = 547
	c                      = 548
	d                      = 549
	e                      = 550
	f                      = 551
	g                      = 552
	h                      = 553
	i                      = 554
	j                      = 555
	k                      = 556
	l                      = 557
	m                      = 558
	n                      = 559
	o                      = 560
	p                      = 561
	q                      = 562
	r                      = 563
	s                      = 564
	t                      = 565
	u                      = 566
	v                      = 567
	w                      = 568
	x                      = 569
	y                      = 570
	z                      = 571
	f1                     = 572
	f2                     = 573
	f3                     = 574
	f4                     = 575
	f5                     = 576
	f6                     = 577
	f7                     = 578
	f8                     = 579
	f9                     = 580
	f10                    = 581
	f11                    = 582
	f12                    = 583
	f13                    = 584
	f14                    = 585
	f15                    = 586
	f16                    = 587
	f17                    = 588
	f18                    = 589
	f19                    = 590
	f20                    = 591
	f21                    = 592
	f22                    = 593
	f23                    = 594
	f24                    = 595
	apostrophe             = 596
	comma                  = 597
	minus                  = 598
	period                 = 599
	slash                  = 600
	semicolon              = 601
	equal                  = 602
	left_bracket           = 603
	backslash              = 604
	right_bracket          = 605
	grave_accent           = 606
	caps_lock              = 607
	scroll_lock            = 608
	num_lock               = 609
	print_screen           = 610
	pause                  = 611
	pad0                   = 612
	pad1                   = 613
	pad2                   = 614
	pad3                   = 615
	pad4                   = 616
	pad5                   = 617
	pad6                   = 618
	pad7                   = 619
	pad8                   = 620
	pad9                   = 621
	pad_decimal            = 622
	pad_divide             = 623
	pad_multiply           = 624
	pad_subtract           = 625
	pad_add                = 626
	pad_enter              = 627
	pad_equal              = 628
	app_back               = 629
	app_forward            = 630
	oem102                 = 631
	gamepad_start          = 632
	gamepad_back           = 633
	gamepad_face_left      = 634
	gamepad_face_right     = 635
	gamepad_face_up        = 636
	gamepad_face_down      = 637
	gamepad_dpad_left      = 638
	gamepad_dpad_right     = 639
	gamepad_dpad_up        = 640
	gamepad_dpad_down      = 641
	gamepad_l1             = 642
	gamepad_r1             = 643
	gamepad_l2             = 644
	gamepad_r2             = 645
	gamepad_l3             = 646
	gamepad_r3             = 647
	gamepad_ls_tick_left   = 648
	gamepad_ls_tick_right  = 649
	gamepad_ls_tick_up     = 650
	gamepad_ls_tick_down   = 651
	gamepad_rs_tick_left   = 652
	gamepad_rs_tick_right  = 653
	gamepad_rs_tick_up     = 654
	gamepad_rs_tick_down   = 655
	mouse_left             = 656
	mouse_right            = 657
	mouse_middle           = 658
	mouse_x1               = 659
	mouse_x2               = 660
	mouse_wheel_x          = 661
	mouse_wheel_y          = 662
	reserved_for_mod_ctrl  = 663
	reserved_for_mod_shift = 664
	reserved_for_mod_alt   = 665
	reserved_for_mod_super = 666
	named_end              = 667
	mod_none               = 0
	mod_ctrl               = 1 << 12
	mod_shift              = 1 << 13
	mod_alt                = 1 << 14
	mod_super              = 1 << 15
	mod_mask_              = 61440
	named_count            = 667 - 512
}

enum InputFlags_ {
	none                    = 0
	repeat                  = 1 << 0
	route_active            = 1 << 10
	route_focused           = 1 << 11
	route_global            = 1 << 12
	route_always            = 1 << 13
	route_over_focused      = 1 << 14
	route_over_active       = 1 << 15
	route_unless_bg_focused = 1 << 16
	route_from_root_window  = 1 << 17
	tooltip                 = 1 << 18
}

enum ConfigFlags_ {
	none                       = 0
	nav_enable_keyboard        = 1 << 0
	nav_enable_gamepad         = 1 << 1
	no_mouse                   = 1 << 4
	no_mouse_cursor_change     = 1 << 5
	no_keyboard                = 1 << 6
	docking_enable             = 1 << 7
	viewports_enable           = 1 << 10
	dpi_enable_scale_viewports = 1 << 14
	dpi_enable_scale_fonts     = 1 << 15
	is_srgb                    = 1 << 20
	is_touch_screen            = 1 << 21
}

enum BackendFlags_ {
	none                       = 0
	has_gamepad                = 1 << 0
	has_mouse_cursors          = 1 << 1
	has_set_mouse_pos          = 1 << 2
	renderer_has_vtx_offset    = 1 << 3
	platform_has_viewports     = 1 << 10
	has_mouse_hovered_viewport = 1 << 11
	renderer_has_viewports     = 1 << 12
}

enum Col_ {
	text
	text_disabled
	window_bg
	child_bg
	popup_bg
	border
	border_shadow
	frame_bg
	frame_bg_hovered
	frame_bg_active
	title_bg
	title_bg_active
	title_bg_collapsed
	menu_bar_bg
	scrollbar_bg
	scrollbar_grab
	scrollbar_grab_hovered
	scrollbar_grab_active
	check_mark
	slider_grab
	slider_grab_active
	button
	button_hovered
	button_active
	header
	header_hovered
	header_active
	separator
	separator_hovered
	separator_active
	resize_grip
	resize_grip_hovered
	resize_grip_active
	tab_hovered
	tab
	tab_selected
	tab_selected_overline
	tab_dimmed
	tab_dimmed_selected
	tab_dimmed_selected_overline
	docking_preview
	docking_empty_bg
	plot_lines
	plot_lines_hovered
	plot_histogram
	plot_histogram_hovered
	table_header_bg
	table_border_strong
	table_border_light
	table_row_bg
	table_row_bg_alt
	text_link
	text_selected_bg
	drag_drop_target
	nav_cursor
	nav_windowing_highlight
	nav_windowing_dim_bg
	modal_window_dim_bg
	count
}

enum StyleVar_ {
	alpha
	disabled_alpha
	window_padding
	window_rounding
	window_border_size
	window_min_size
	window_title_align
	child_rounding
	child_border_size
	popup_rounding
	popup_border_size
	frame_padding
	frame_rounding
	frame_border_size
	item_spacing
	item_inner_spacing
	indent_spacing
	cell_padding
	scrollbar_size
	scrollbar_rounding
	grab_min_size
	grab_rounding
	image_border_size
	tab_rounding
	tab_border_size
	tab_bar_border_size
	tab_bar_overline_size
	table_angled_headers_angle
	table_angled_headers_text_align
	button_text_align
	selectable_text_align
	separator_text_border_size
	separator_text_align
	separator_text_padding
	docking_separator_size
	count
}

enum ButtonFlags_ {
	none                = 0
	mouse_button_left   = 1 << 0
	mouse_button_right  = 1 << 1
	mouse_button_middle = 1 << 2
	mouse_button_mask_  = 1 << 0 | 1 << 1 | 1 << 2
	enable_nav          = 1 << 3
}

enum ColorEditFlags_ {
	none               = 0
	no_alpha           = 1 << 1
	no_picker          = 1 << 2
	no_options         = 1 << 3
	no_small_preview   = 1 << 4
	no_inputs          = 1 << 5
	no_tooltip         = 1 << 6
	no_label           = 1 << 7
	no_side_preview    = 1 << 8
	no_drag_drop       = 1 << 9
	no_border          = 1 << 10
	alpha_opaque       = 1 << 11
	alpha_no_bg        = 1 << 12
	alpha_preview_half = 1 << 13
	alpha_bar          = 1 << 16
	hdr                = 1 << 19
	display_rgb        = 1 << 20
	display_hsv        = 1 << 21
	display_hex        = 1 << 22
	uint8              = 1 << 23
	float              = 1 << 24
	picker_hue_bar     = 1 << 25
	picker_hue_wheel   = 1 << 26
	input_rgb          = 1 << 27
	input_hsv          = 1 << 28
	default_options_   = 1 << 23 | 1 << 20 | 1 << 27 | 1 << 25
	alpha_mask_        = 1 << 1 | 1 << 11 | 1 << 12 | 1 << 13
	display_mask_      = 1 << 20 | 1 << 21 | 1 << 22
	data_type_mask_    = 1 << 23 | 1 << 24
	picker_mask_       = 1 << 26 | 1 << 25
	input_mask_        = 1 << 27 | 1 << 28
}

enum SliderFlags_ {
	none               = 0
	logarithmic        = 1 << 5
	no_round_to_format = 1 << 6
	no_input           = 1 << 7
	wrap_around        = 1 << 8
	clamp_on_input     = 1 << 9
	clamp_zero_range   = 1 << 10
	no_speed_tweaks    = 1 << 11
	always_clamp       = 1 << 9 | 1 << 10
	invalid_mask_      = 1879048207
}

enum MouseButton_ {
	left   = 0
	right  = 1
	middle = 2
	count  = 5
}

enum MouseCursor_ {
	none  = -1
	arrow = 0
	text_input
	resize_all
	resize_ns
	resize_ew
	resize_nesw
	resize_nwse
	hand
	wait
	progress
	not_allowed
	count
}

enum MouseSource {
	mouse        = 0
	touch_screen = 1
	pen          = 2
	count        = 3
}

enum Cond_ {
	none           = 0
	always         = 1 << 0
	once           = 1 << 1
	first_use_ever = 1 << 2
	appearing      = 1 << 3
}

enum TableFlags_ {
	none                            = 0
	resizable                       = 1 << 0
	reorderable                     = 1 << 1
	hideable                        = 1 << 2
	sortable                        = 1 << 3
	no_saved_settings               = 1 << 4
	context_menu_in_body            = 1 << 5
	row_bg                          = 1 << 6
	borders_inner_h                 = 1 << 7
	borders_outer_h                 = 1 << 8
	borders_inner_v                 = 1 << 9
	borders_outer_v                 = 1 << 10
	borders_h                       = 1 << 7 | 1 << 8
	borders_v                       = 1 << 9 | 1 << 10
	borders_inner                   = 1 << 9 | 1 << 7
	borders_outer                   = 1 << 10 | 1 << 8
	borders                         = 1 << 9 | 1 << 7 | 1 << 10 | 1 << 8
	no_borders_in_body              = 1 << 11
	no_borders_in_body_until_resize = 1 << 12
	sizing_fixed_fit                = 1 << 13
	sizing_fixed_same               = 2 << 13
	sizing_stretch_prop             = 3 << 13
	sizing_stretch_same             = 4 << 13
	no_host_extend_x                = 1 << 16
	no_host_extend_y                = 1 << 17
	no_keep_columns_visible         = 1 << 18
	precise_widths                  = 1 << 19
	no_clip                         = 1 << 20
	pad_outer_x                     = 1 << 21
	no_pad_outer_x                  = 1 << 22
	no_pad_inner_x                  = 1 << 23
	scroll_x                        = 1 << 24
	scroll_y                        = 1 << 25
	sort_multi                      = 1 << 26
	sort_tristate                   = 1 << 27
	highlight_hovered_column        = 1 << 28
	sizing_mask_                    = 1 << 13 | 2 << 13 | 3 << 13 | 4 << 13
}

enum TableColumnFlags_ {
	none                   = 0
	disabled               = 1 << 0
	default_hide           = 1 << 1
	default_sort           = 1 << 2
	width_stretch          = 1 << 3
	width_fixed            = 1 << 4
	no_resize              = 1 << 5
	no_reorder             = 1 << 6
	no_hide                = 1 << 7
	no_clip                = 1 << 8
	no_sort                = 1 << 9
	no_sort_ascending      = 1 << 10
	no_sort_descending     = 1 << 11
	no_header_label        = 1 << 12
	no_header_width        = 1 << 13
	prefer_sort_ascending  = 1 << 14
	prefer_sort_descending = 1 << 15
	indent_enable          = 1 << 16
	indent_disable         = 1 << 17
	angled_header          = 1 << 18
	is_enabled             = 1 << 24
	is_visible             = 1 << 25
	is_sorted              = 1 << 26
	is_hovered             = 1 << 27
	width_mask_            = 1 << 3 | 1 << 4
	indent_mask_           = 1 << 16 | 1 << 17
	status_mask_           = 1 << 24 | 1 << 25 | 1 << 26 | 1 << 27
	no_direct_resize_      = 1 << 30
}

enum TableRowFlags_ {
	none    = 0
	headers = 1 << 0
}

enum TableBgTarget_ {
	none    = 0
	row_bg0 = 1
	row_bg1 = 2
	cell_bg = 3
}

struct TableSortSpecs {
	specs      &TableColumnSortSpecs
	specsCount int
	specsDirty bool
}

struct TableColumnSortSpecs {
	columnUserID  ID
	columnIndex   ImS16
	sortOrder     ImS16
	sortDirection SortDirection
}

struct Style {
	alpha                            f32
	disabledAlpha                    f32
	windowPadding                    ImVec2
	windowRounding                   f32
	windowBorderSize                 f32
	windowBorderHoverPadding         f32
	windowMinSize                    ImVec2
	windowTitleAlign                 ImVec2
	windowMenuButtonPosition         Dir
	childRounding                    f32
	childBorderSize                  f32
	popupRounding                    f32
	popupBorderSize                  f32
	framePadding                     ImVec2
	frameRounding                    f32
	frameBorderSize                  f32
	itemSpacing                      ImVec2
	itemInnerSpacing                 ImVec2
	cellPadding                      ImVec2
	touchExtraPadding                ImVec2
	indentSpacing                    f32
	columnsMinSpacing                f32
	scrollbarSize                    f32
	scrollbarRounding                f32
	grabMinSize                      f32
	grabRounding                     f32
	logSliderDeadzone                f32
	imageBorderSize                  f32
	tabRounding                      f32
	tabBorderSize                    f32
	tabCloseButtonMinWidthSelected   f32
	tabCloseButtonMinWidthUnselected f32
	tabBarBorderSize                 f32
	tabBarOverlineSize               f32
	tableAngledHeadersAngle          f32
	tableAngledHeadersTextAlign      ImVec2
	colorButtonPosition              Dir
	buttonTextAlign                  ImVec2
	selectableTextAlign              ImVec2
	separatorTextBorderSize          f32
	separatorTextAlign               ImVec2
	separatorTextPadding             ImVec2
	displayWindowPadding             ImVec2
	displaySafeAreaPadding           ImVec2
	dockingSeparatorSize             f32
	mouseCursorScale                 f32
	antiAliasedLines                 bool
	antiAliasedLinesUseTex           bool
	antiAliasedFill                  bool
	curveTessellationTol             f32
	circleTessellationMaxError       f32
	colors                           [58]C.ImVec4
	hoverStationaryDelay             f32
	hoverDelayShort                  f32
	hoverDelayNormal                 f32
	hoverFlagsForTooltipMouse        HoveredFlags
	hoverFlagsForTooltipNav          HoveredFlags
}

struct KeyData {
	down             bool
	downDuration     f32
	downDurationPrev f32
	analogValue      f32
}

struct ImVector_ImWchar {
	size     int
	capacity int
	data     &C.ImWchar
}

struct IO {
	configFlags                                   ConfigFlags
	backendFlags                                  BackendFlags
	displaySize                                   ImVec2
	deltaTime                                     f32
	iniSavingRate                                 f32
	iniFilename                                   &i8
	logFilename                                   &i8
	userData                                      voidptr
	fonts                                         &ImFontAtlas
	fontGlobalScale                               f32
	fontAllowUserScaling                          bool
	fontDefault                                   &ImFont
	displayFramebufferScale                       ImVec2
	configNavSwapGamepadButtons                   bool
	configNavMoveSetMousePos                      bool
	configNavCaptureKeyboard                      bool
	configNavEscapeClearFocusItem                 bool
	configNavEscapeClearFocusWindow               bool
	configNavCursorVisibleAuto                    bool
	configNavCursorVisibleAlways                  bool
	configDockingNoSplit                          bool
	configDockingWithShift                        bool
	configDockingAlwaysTabBar                     bool
	configDockingTransparentPayload               bool
	configViewportsNoAutoMerge                    bool
	configViewportsNoTaskBarIcon                  bool
	configViewportsNoDecoration                   bool
	configViewportsNoDefaultParent                bool
	mouseDrawCursor                               bool
	configMacOSXBehaviors                         bool
	configInputTrickleEventQueue                  bool
	configInputTextCursorBlink                    bool
	configInputTextEnterKeepActive                bool
	configDragClickToInputText                    bool
	configWindowsResizeFromEdges                  bool
	configWindowsMoveFromTitleBarOnly             bool
	configWindowsCopyContentsWithCtrlC            bool
	configScrollbarScrollByPage                   bool
	configMemoryCompactTimer                      f32
	mouseDoubleClickTime                          f32
	mouseDoubleClickMaxDist                       f32
	mouseDragThreshold                            f32
	keyRepeatDelay                                f32
	keyRepeatRate                                 f32
	configErrorRecovery                           bool
	configErrorRecoveryEnableAssert               bool
	configErrorRecoveryEnableDebugLog             bool
	configErrorRecoveryEnableTooltip              bool
	configDebugIsDebuggerPresent                  bool
	configDebugHighlightIdConflicts               bool
	configDebugHighlightIdConflictsShowItemPicker bool
	configDebugBeginReturnValueOnce               bool
	configDebugBeginReturnValueLoop               bool
	configDebugIgnoreFocusLoss                    bool
	configDebugIniSettings                        bool
	backendPlatformName                           &i8
	backendRendererName                           &i8
	backendPlatformUserData                       voidptr
	backendRendererUserData                       voidptr
	backendLanguageUserData                       voidptr
	wantCaptureMouse                              bool
	wantCaptureKeyboard                           bool
	wantTextInput                                 bool
	wantSetMousePos                               bool
	wantSaveIniSettings                           bool
	navActive                                     bool
	navVisible                                    bool
	framerate                                     f32
	metricsRenderVertices                         int
	metricsRenderIndices                          int
	metricsRenderWindows                          int
	metricsActiveWindows                          int
	mouseDelta                                    ImVec2
	ctx                                           &Context
	mousePos                                      ImVec2
	mouseDown                                     [5]bool
	mouseWheel                                    f32
	mouseWheelH                                   f32
	mouseSource                                   MouseSource
	mouseHoveredViewport                          ID
	keyCtrl                                       bool
	keyShift                                      bool
	keyAlt                                        bool
	keySuper                                      bool
	keyMods                                       KeyChord
	keysData                                      [155]KeyData
	wantCaptureMouseUnlessPopupClose              bool
	mousePosPrev                                  ImVec2
	mouseClickedPos                               [5]ImVec2
	mouseClickedTime                              [5]f64
	mouseClicked                                  [5]bool
	mouseDoubleClicked                            [5]bool
	mouseClickedCount                             [5]ImU16
	mouseClickedLastCount                         [5]ImU16
	mouseReleased                                 [5]bool
	mouseReleasedTime                             [5]f64
	mouseDownOwned                                [5]bool
	mouseDownOwnedUnlessPopupClose                [5]bool
	mouseWheelRequestAxisSwap                     bool
	mouseCtrlLeftAsRightClick                     bool
	mouseDownDuration                             [5]f32
	mouseDownDurationPrev                         [5]f32
	mouseDragMaxDistanceAbs                       [5]ImVec2
	mouseDragMaxDistanceSqr                       [5]f32
	penPressure                                   f32
	appFocusLost                                  bool
	appAcceptingEvents                            bool
	inputQueueSurrogate                           ImWchar16
	inputQueueCharacters                          ImVector_ImWchar
}

struct ImGuiInputTextCallbackData {
	ctx            &Context
	eventFlag      InputTextFlags
	flags          InputTextFlags
	userData       voidptr
	eventChar      C.ImWchar
	eventKey       Key
	buf            &i8
	bufTextLen     int
	bufSize        int
	bufDirty       bool
	cursorPos      int
	selectionStart int
	selectionEnd   int
}

struct ImGuiSizeCallbackData {
	userData    voidptr
	pos         ImVec2
	currentSize ImVec2
	desiredSize ImVec2
}

struct WindowClass {
	classId                    ID
	parentViewportId           ID
	focusRouteParentWindowId   ID
	viewportFlagsOverrideSet   ViewportFlags
	viewportFlagsOverrideClear ViewportFlags
	tabItemFlagsOverrideSet    TabItemFlags
	dockNodeFlagsOverrideSet   DockNodeFlags
	dockingAlwaysTabBar        bool
	dockingAllowUnclassed      bool
}

struct Payload {
	data           voidptr
	dataSize       int
	sourceId       ID
	sourceParentId ID
	dataFrameCount int
	dataType       [33]i8
	preview        bool
	delivery       bool
}

struct OnceUponAFrame {
	refFrame int
}

struct TextRange {
	b &i8
	e &i8
}

struct ImVector_ImGuiTextRange {
	size     int
	capacity int
	data     &TextRange
}

struct ImVector_char {
	size     int
	capacity int
	data     &i8
}

struct TextBuffer {
	buf ImVector_char
}

struct StoragePair {
	key ID
}

struct ImVector_ImGuiStoragePair {
	size     int
	capacity int
	data     &StoragePair
}

struct Storage {
	data ImVector_ImGuiStoragePair
}

struct ListClipper {
	ctx              &Context
	displayStart     int
	displayEnd       int
	itemsCount       int
	itemsHeight      f32
	startPosY        f32
	startSeekOffsetY f64
	tempData         voidptr
}

struct ImColor {
	value C.ImVec4
}

enum MultiSelectFlags_ {
	none                      = 0
	single_select             = 1 << 0
	no_select_all             = 1 << 1
	no_range_select           = 1 << 2
	no_auto_select            = 1 << 3
	no_auto_clear             = 1 << 4
	no_auto_clear_on_reselect = 1 << 5
	box_select1d              = 1 << 6
	box_select2d              = 1 << 7
	box_select_no_scroll      = 1 << 8
	clear_on_escape           = 1 << 9
	clear_on_click_void       = 1 << 10
	scope_window              = 1 << 11
	scope_rect                = 1 << 12
	select_on_click           = 1 << 13
	select_on_click_release   = 1 << 14
	nav_wrap_x                = 1 << 16
}

struct ImVector_ImGuiSelectionRequest {
	size     int
	capacity int
	data     &SelectionRequest
}

struct MultiSelectIO {
	requests      ImVector_ImGuiSelectionRequest
	rangeSrcItem  SelectionUserData
	navIdItem     SelectionUserData
	navIdSelected bool
	rangeSrcReset bool
	itemsCount    int
}

enum SelectionRequestType {
	none = 0
	set_all
	set_range
}

struct SelectionRequest {
	type           SelectionRequestType
	selected       bool
	rangeDirection ImS8
	rangeFirstItem SelectionUserData
	rangeLastItem  SelectionUserData
}

struct SelectionBasicStorage {
	size                    int
	preserveOrder           bool
	userData                voidptr
	adapterIndexToStorageId fn (&SelectionBasicStorage, int) ID
	_SelectionOrder         int
	_Storage                Storage
}

struct ImDrawIdx {
	userData               voidptr
	adapterSetItemSelected fn (&C.ImGuiSelectionExternalStorage, int, bool)
}

type ImDrawCallback = fn (&ImDrawList, &ImDrawCmd)

struct ImDrawCmd {
	clipRect               C.ImVec4
	textureId              ImTextureID
	vtxOffset              u32
	idxOffset              u32
	elemCount              u32
	userCallback           ImDrawCallback
	userCallbackData       voidptr
	userCallbackDataSize   int
	userCallbackDataOffset int
}

struct ImDrawVert {
	pos ImVec2
	uv  ImVec2
	col ImU32
}

struct ImDrawCmdHeader {
	clipRect  C.ImVec4
	textureId ImTextureID
	vtxOffset u32
}

struct ImVector_ImDrawCmd {
	size     int
	capacity int
	data     &ImDrawCmd
}

struct ImVector_ImDrawIdx {
	size     int
	capacity int
	data     &ImDrawIdx
}

struct ImDrawChannel {
	_CmdBuffer ImVector_ImDrawCmd
	_IdxBuffer ImVector_ImDrawIdx
}

struct ImVector_ImDrawChannel {
	size     int
	capacity int
	data     &ImDrawChannel
}

struct ImDrawListSplitter {
	_Current  int
	_Count    int
	_Channels ImVector_ImDrawChannel
}

enum ImDrawFlags_ {
	none                       = 0
	closed                     = 1 << 0
	round_corners_top_left     = 1 << 4
	round_corners_top_right    = 1 << 5
	round_corners_bottom_left  = 1 << 6
	round_corners_bottom_right = 1 << 7
	round_corners_none         = 1 << 8
	round_corners_top          = 1 << 4 | 1 << 5
	round_corners_bottom       = 1 << 6 | 1 << 7
	round_corners_left         = 1 << 6 | 1 << 4
	round_corners_right        = 1 << 7 | 1 << 5
	round_corners_all          = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	round_corners_default_     = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	round_corners_mask_        = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8
}

enum ImDrawListFlags_ {
	none                       = 0
	anti_aliased_lines         = 1 << 0
	anti_aliased_lines_use_tex = 1 << 1
	anti_aliased_fill          = 1 << 2
	allow_vtx_offset           = 1 << 3
}

struct ImVector_ImDrawVert {
	size     int
	capacity int
	data     &ImDrawVert
}

struct ImVector_ImVec2 {
	size     int
	capacity int
	data     &ImVec2
}

struct ImVector_ImVec4 {
	size     int
	capacity int
	data     &C.ImVec4
}

struct ImVector_ImTextureID {
	size     int
	capacity int
	data     &ImTextureID
}

struct ImVector_ImU8 {
	size     int
	capacity int
	data     &ImU8
}

struct ImDrawList {
	cmdBuffer         ImVector_ImDrawCmd
	idxBuffer         ImVector_ImDrawIdx
	vtxBuffer         ImVector_ImDrawVert
	flags             ImDrawListFlags
	_VtxCurrentIdx    u32
	_Data             &ImDrawListSharedData
	_VtxWritePtr      &ImDrawVert
	_IdxWritePtr      &ImDrawIdx
	_Path             ImVector_ImVec2
	_CmdHeader        ImDrawCmdHeader
	_Splitter         ImDrawListSplitter
	_ClipRectStack    ImVector_ImVec4
	_TextureIdStack   ImVector_ImTextureID
	_CallbacksDataBuf ImVector_ImU8
	_FringeScale      f32
	_OwnerName        &i8
}

struct ImVector_ImDrawListPtr {
	size     int
	capacity int
	data     &&ImDrawList
}

struct ImDrawData {
	valid            bool
	cmdListsCount    int
	totalIdxCount    int
	totalVtxCount    int
	cmdLists         ImVector_ImDrawListPtr
	displayPos       ImVec2
	displaySize      ImVec2
	framebufferScale ImVec2
	ownerViewport    &Viewport
}

struct ImFontConfig {
	fontData             voidptr
	fontDataSize         int
	fontDataOwnedByAtlas bool
	mergeMode            bool
	pixelSnapH           bool
	fontNo               int
	oversampleH          int
	oversampleV          int
	sizePixels           f32
	glyphOffset          ImVec2
	glyphRanges          &C.ImWchar
	glyphMinAdvanceX     f32
	glyphMaxAdvanceX     f32
	glyphExtraAdvanceX   f32
	fontBuilderFlags     u32
	rasterizerMultiply   f32
	rasterizerDensity    f32
	ellipsisChar         C.ImWchar
	name                 [40]i8
	dstFont              &ImFont
}

struct ImFontGlyph {
	colored   u32
	visible   u32
	codepoint u32
	advanceX  f32
	x0        f32
	y0        f32
	x1        f32
	y1        f32
	u0        f32
	v0        f32
	u1        f32
	v1        f32
}

struct ImVector_ImU32 {
	size     int
	capacity int
	data     &ImU32
}

struct ImFontGlyphRangesBuilder {
	usedChars ImVector_ImU32
}

struct ImFontAtlasCustomRect {
	x             u16
	y             u16
	width         u16
	height        u16
	glyphID       u32
	glyphColored  u32
	glyphAdvanceX f32
	glyphOffset   ImVec2
	font          &ImFont
}

enum ImFontAtlasFlags_ {
	none                   = 0
	no_power_of_two_height = 1 << 0
	no_mouse_cursors       = 1 << 1
	no_baked_lines         = 1 << 2
}

struct ImVector_ImFontPtr {
	size     int
	capacity int
	data     &&ImFont
}

struct ImVector_ImFontAtlasCustomRect {
	size     int
	capacity int
	data     &ImFontAtlasCustomRect
}

struct ImVector_ImFontConfig {
	size     int
	capacity int
	data     &ImFontConfig
}

struct ImFontAtlas {
	flags              ImFontAtlasFlags
	texID              ImTextureID
	texDesiredWidth    int
	texGlyphPadding    int
	userData           voidptr
	locked             bool
	texReady           bool
	texPixelsUseColors bool
	texPixelsAlpha8    &u8
	texPixelsRGBA32    &u32
	texWidth           int
	texHeight          int
	texUvScale         ImVec2
	texUvWhitePixel    ImVec2
	fonts              ImVector_ImFontPtr
	customRects        ImVector_ImFontAtlasCustomRect
	sources            ImVector_ImFontConfig
	texUvLines         [33]C.ImVec4
	fontBuilderIO      &ImFontBuilderIO
	fontBuilderFlags   u32
	packIdMouseCursors int
	packIdLines        int
}

struct ImVector_float {
	size     int
	capacity int
	data     &f32
}

struct ImVector_ImU16 {
	size     int
	capacity int
	data     &ImU16
}

struct ImVector_ImFontGlyph {
	size     int
	capacity int
	data     &ImFontGlyph
}

struct ImFont {
	indexAdvanceX       ImVector_float
	fallbackAdvanceX    f32
	fontSize            f32
	indexLookup         ImVector_ImU16
	glyphs              ImVector_ImFontGlyph
	fallbackGlyph       &ImFontGlyph
	containerAtlas      &ImFontAtlas
	sources             &ImFontConfig
	sourcesCount        i16
	ellipsisCharCount   i16
	ellipsisChar        C.ImWchar
	fallbackChar        C.ImWchar
	ellipsisWidth       f32
	ellipsisCharStep    f32
	scale               f32
	ascent              f32
	descent             f32
	metricsTotalSurface int
	dirtyLookupTables   bool
	used8kPagesMap      [17]ImU8
}

enum ViewportFlags_ {
	none                   = 0
	is_platform_window     = 1 << 0
	is_platform_monitor    = 1 << 1
	owned_by_app           = 1 << 2
	no_decoration          = 1 << 3
	no_task_bar_icon       = 1 << 4
	no_focus_on_appearing  = 1 << 5
	no_focus_on_click      = 1 << 6
	no_inputs              = 1 << 7
	no_renderer_clear      = 1 << 8
	no_auto_merge          = 1 << 9
	top_most               = 1 << 10
	can_host_other_windows = 1 << 11
	is_minimized           = 1 << 12
	is_focused             = 1 << 13
}

struct Viewport {
	iD                    ID
	flags                 ViewportFlags
	pos                   ImVec2
	size                  ImVec2
	workPos               ImVec2
	workSize              ImVec2
	dpiScale              f32
	parentViewportId      ID
	drawData              &ImDrawData
	rendererUserData      voidptr
	platformUserData      voidptr
	platformHandle        voidptr
	platformHandleRaw     voidptr
	platformWindowCreated bool
	platformRequestMove   bool
	platformRequestResize bool
	platformRequestClose  bool
}

struct ImVector_ImGuiPlatformMonitor {
	size     int
	capacity int
	data     &PlatformMonitor
}

struct ImVector_ImGuiViewportPtr {
	size     int
	capacity int
	data     &&Viewport
}

struct PlatformIO {
	platform_GetClipboardTextFn      fn (&Context) &i8
	platform_SetClipboardTextFn      fn (&Context, &i8)
	platform_ClipboardUserData       voidptr
	platform_OpenInShellFn           fn (&Context, &i8) bool
	platform_OpenInShellUserData     voidptr
	platform_SetImeDataFn            fn (&Context, &Viewport, &PlatformImeData)
	platform_ImeUserData             voidptr
	platform_LocaleDecimalPoint      C.ImWchar
	renderer_RenderState             voidptr
	platform_CreateWindow            fn (&Viewport)
	platform_DestroyWindow           fn (&Viewport)
	platform_ShowWindow              fn (&Viewport)
	platform_SetWindowPos            fn (&Viewport, ImVec2)
	platform_GetWindowPos            fn (&Viewport) ImVec2
	platform_SetWindowSize           fn (&Viewport, ImVec2)
	platform_GetWindowSize           fn (&Viewport) ImVec2
	platform_SetWindowFocus          fn (&Viewport)
	platform_GetWindowFocus          fn (&Viewport) bool
	platform_GetWindowMinimized      fn (&Viewport) bool
	platform_SetWindowTitle          fn (&Viewport, &i8)
	platform_SetWindowAlpha          fn (&Viewport, f32)
	platform_UpdateWindow            fn (&Viewport)
	platform_RenderWindow            fn (&Viewport, voidptr)
	platform_SwapBuffers             fn (&Viewport, voidptr)
	platform_GetWindowDpiScale       fn (&Viewport) f32
	platform_OnChangedViewport       fn (&Viewport)
	platform_GetWindowWorkAreaInsets fn (&Viewport) C.ImVec4
	platform_CreateVkSurface         fn (&Viewport, ImU64, voidptr, &ImU64) int
	renderer_CreateWindow            fn (&Viewport)
	renderer_DestroyWindow           fn (&Viewport)
	renderer_SetWindowSize           fn (&Viewport, ImVec2)
	renderer_RenderWindow            fn (&Viewport, voidptr)
	renderer_SwapBuffers             fn (&Viewport, voidptr)
	monitors                         ImVector_ImGuiPlatformMonitor
	viewports                        ImVector_ImGuiViewportPtr
}

struct PlatformMonitor {
	mainPos        ImVec2
	mainSize       ImVec2
	workPos        ImVec2
	workSize       ImVec2
	dpiScale       f32
	platformHandle voidptr
}

struct PlatformImeData {
	wantVisible     bool
	inputPos        ImVec2
	inputLineHeight f32
}

type DataAuthority = int
type LayoutType = int
type ActivateFlags = int
type DebugLogFlags = int
type FocusRequestFlags = int
type ItemStatusFlags = int
type OldColumnFlags = int
type LogFlags = int
type NavRenderCursorFlags = int
type NavMoveFlags = int
type NextItemDataFlags = int
type NextWindowDataFlags = int
type ScrollFlags = int
type SeparatorFlags = int
type TextFlags = int
type TooltipFlags = int
type TypingSelectFlags = int
type WindowRefreshFlags = int

@[weak]
__global GImGui &Context

type ImFileHandle = &C.FILE

struct ImVec1 {
	x f32
}

struct ImVec2ih {
	x i16
	y i16
}

struct ImBitArrayPtr {
	min ImVec2
	max ImVec2
}

struct ImPoolIdx {
	storage ImVector_ImU32
}

struct ImVector_int {
	size     int
	capacity int
	data     &int
}

struct TextIndex {
	lineOffsets ImVector_int
	endOffset   int
}

struct ImDrawListSharedData {
	texUvWhitePixel       ImVec2
	texUvLines            &C.ImVec4
	font                  &ImFont
	fontSize              f32
	fontScale             f32
	curveTessellationTol  f32
	circleSegmentMaxError f32
	initialFringeScale    f32
	initialFlags          ImDrawListFlags
	clipRectFullscreen    C.ImVec4
	tempBuffer            ImVector_ImVec2
	arcFastVtx            [48]ImVec2
	arcFastRadiusCutoff   f32
	circleSegmentCounts   [64]ImU8
}

struct ImDrawDataBuilder {
	layers     [2]&ImVector_ImDrawListPtr
	layerData1 ImVector_ImDrawListPtr
}

struct StyleVarInfo {
	count    ImU32
	dataType DataType
	offset   ImU32
}

struct ColorMod {
	col         Col
	backupValue C.ImVec4
}

struct StyleMod {
	varIdx StyleVar
}

struct DataTypeStorage {
	data [8]ImU8
}

struct DataTypeInfo {
	size     usize
	name     &i8
	printFmt &i8
	scanFmt  &i8
}

enum DataTypePrivate_ {
	pointer = int(DataType_.count)
	id
}

enum ItemFlagsPrivate_ {
	disabled                   = 1 << 10
	read_only                  = 1 << 11
	mixed_value                = 1 << 12
	no_window_hoverable_check  = 1 << 13
	allow_overlap              = 1 << 14
	no_nav_disable_mouse_hover = 1 << 15
	no_mark_edited             = 1 << 16
	inputable                  = 1 << 20
	has_selection_user_data    = 1 << 21
	is_multi_select            = 1 << 22
	default_                   = 1 << 4
}

enum ItemStatusFlags_ {
	none              = 0
	hovered_rect      = 1 << 0
	has_display_rect  = 1 << 1
	edited            = 1 << 2
	toggled_selection = 1 << 3
	toggled_open      = 1 << 4
	has_deactivated   = 1 << 5
	deactivated       = 1 << 6
	hovered_window    = 1 << 7
	visible           = 1 << 8
	has_clip_rect     = 1 << 9
	has_shortcut      = 1 << 10
}

enum HoveredFlagsPrivate_ {
	delay_mask_                        = 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
	allowed_mask_for_is_window_hovered = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 7 | 1 << 12 | 1 << 13
	allowed_mask_for_is_item_hovered   = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
}

enum InputTextFlagsPrivate_ {
	multiline              = 1 << 26
	merged_item            = 1 << 27
	localize_decimal_point = 1 << 28
}

enum ButtonFlagsPrivate_ {
	pressed_on_click                  = 1 << 4
	pressed_on_click_release          = 1 << 5
	pressed_on_click_release_anywhere = 1 << 6
	pressed_on_release                = 1 << 7
	pressed_on_double_click           = 1 << 8
	pressed_on_drag_drop_hold         = 1 << 9
	flatten_children                  = 1 << 11
	allow_overlap                     = 1 << 12
	align_text_base_line              = 1 << 15
	no_key_mods_allowed               = 1 << 16
	no_holding_active_id              = 1 << 17
	no_nav_focus                      = 1 << 18
	no_hovered_on_focus               = 1 << 19
	no_set_key_owner                  = 1 << 20
	no_test_key_owner                 = 1 << 21
	pressed_on_mask_                  = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8 | 1 << 9
	pressed_on_default_               = 1 << 5
}

enum ComboFlagsPrivate_ {
	custom_preview = 1 << 20
}

enum SliderFlagsPrivate_ {
	vertical  = 1 << 20
	read_only = 1 << 21
}

enum SelectableFlagsPrivate_ {
	no_holding_active_id     = 1 << 20
	select_on_nav            = 1 << 21
	select_on_click          = 1 << 22
	select_on_release        = 1 << 23
	span_avail_width         = 1 << 24
	set_nav_id_on_hover      = 1 << 25
	no_pad_with_half_spacing = 1 << 26
	no_set_key_owner         = 1 << 27
}

enum TreeNodeFlagsPrivate_ {
	clip_label_for_trailing_button = 1 << 28
	upside_down_arrow              = 1 << 29
	open_on_mask_                  = 1 << 6 | 1 << 7
}

enum SeparatorFlags_ {
	none             = 0
	horizontal       = 1 << 0
	vertical         = 1 << 1
	span_all_columns = 1 << 2
}

enum FocusRequestFlags_ {
	none                  = 0
	restore_focused_child = 1 << 0
	unless_below_modal    = 1 << 1
}

enum TextFlags_ {
	none                            = 0
	no_width_for_large_clipped_text = 1 << 0
}

enum TooltipFlags_ {
	none              = 0
	override_previous = 1 << 1
}

enum LayoutType_ {
	horizontal = 0
	vertical   = 1
}

enum LogFlags_ {
	none             = 0
	output_tty       = 1 << 0
	output_file      = 1 << 1
	output_buffer    = 1 << 2
	output_clipboard = 1 << 3
	output_mask_     = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
}

enum Axis {
	none = -1
	x    = 0
	y    = 1
}

enum PlotType {
	lines
	histogram
}

struct ComboPreviewData {
	previewRect                  C.ImRect
	backupCursorPos              ImVec2
	backupCursorMaxPos           ImVec2
	backupCursorPosPrevLine      ImVec2
	backupPrevLineTextBaseOffset f32
	backupLayout                 LayoutType
}

struct GroupData {
	windowID                     ID
	backupCursorPos              ImVec2
	backupCursorMaxPos           ImVec2
	backupCursorPosPrevLine      ImVec2
	backupIndent                 ImVec1
	backupGroupOffset            ImVec1
	backupCurrLineSize           ImVec2
	backupCurrLineTextBaseOffset f32
	backupActiveIdIsAlive        ID
	backupDeactivatedIdIsAlive   bool
	backupHoveredIdIsAlive       bool
	backupIsSameLine             bool
	emitItem                     bool
}

struct MenuColumns {
	totalWidth     ImU32
	nextTotalWidth ImU32
	spacing        ImU16
	offsetIcon     ImU16
	offsetLabel    ImU16
	offsetShortcut ImU16
	offsetMark     ImU16
	widths         [4]ImU16
}

struct InputTextDeactivatedState {
	iD    ID
	textA ImVector_char
}

type ImStbTexteditState = voidptr

struct InputTextState {
	ctx                  &Context
	stb                  &ImStbTexteditState
	flags                InputTextFlags
	iD                   ID
	textLen              int
	textSrc              &i8
	textA                ImVector_char
	textToRevertTo       ImVector_char
	callbackTextBackup   ImVector_char
	bufCapacity          int
	scroll               ImVec2
	cursorAnim           f32
	cursorFollow         bool
	selectedAllMouseLock bool
	edited               bool
	wantReloadUserBuf    bool
	reloadSelectionStart int
	reloadSelectionEnd   int
}

enum WindowRefreshFlags_ {
	none                 = 0
	try_to_avoid_refresh = 1 << 0
	refresh_on_hover     = 1 << 1
	refresh_on_focus     = 1 << 2
}

enum NextWindowDataFlags_ {
	none                = 0
	has_pos             = 1 << 0
	has_size            = 1 << 1
	has_content_size    = 1 << 2
	has_collapsed       = 1 << 3
	has_size_constraint = 1 << 4
	has_focus           = 1 << 5
	has_bg_alpha        = 1 << 6
	has_scroll          = 1 << 7
	has_window_flags    = 1 << 8
	has_child_flags     = 1 << 9
	has_refresh_policy  = 1 << 10
	has_viewport        = 1 << 11
	has_dock            = 1 << 12
	has_window_class    = 1 << 13
}

struct NextWindowData {
	hasFlags             NextWindowDataFlags
	posCond              Cond
	sizeCond             Cond
	collapsedCond        Cond
	dockCond             Cond
	posVal               ImVec2
	posPivotVal          ImVec2
	sizeVal              ImVec2
	contentSizeVal       ImVec2
	scrollVal            ImVec2
	windowFlags          WindowFlags
	childFlags           ChildFlags
	posUndock            bool
	collapsedVal         bool
	sizeConstraintRect   C.ImRect
	sizeCallback         C.ImGuiSizeCallback
	sizeCallbackUserData voidptr
	bgAlphaVal           f32
	viewportId           ID
	dockId               ID
	windowClass          WindowClass
	menuBarOffsetMinVal  ImVec2
	refreshFlagsVal      WindowRefreshFlags
}

enum NextItemDataFlags_ {
	none           = 0
	has_width      = 1 << 0
	has_open       = 1 << 1
	has_shortcut   = 1 << 2
	has_ref_val    = 1 << 3
	has_storage_id = 1 << 4
}

struct NextItemData {
	hasFlags          NextItemDataFlags
	itemFlags         ItemFlags
	focusScopeId      ID
	selectionUserData SelectionUserData
	width             f32
	shortcut          KeyChord
	shortcutFlags     InputFlags
	openVal           bool
	openCond          ImU8
	refVal            DataTypeStorage
	storageId         ID
}

struct LastItemData {
	iD          ID
	itemFlags   ItemFlags
	statusFlags ItemStatusFlags
	rect        C.ImRect
	navRect     C.ImRect
	displayRect C.ImRect
	clipRect    C.ImRect
	shortcut    KeyChord
}

struct TreeNodeStackData {
	iD        ID
	treeFlags TreeNodeFlags
	itemFlags ItemFlags
	navRect   C.ImRect
}

struct ErrorRecoveryState {
	sizeOfWindowStack     i16
	sizeOfIDStack         i16
	sizeOfTreeStack       i16
	sizeOfColorStack      i16
	sizeOfStyleVarStack   i16
	sizeOfFontStack       i16
	sizeOfFocusScopeStack i16
	sizeOfGroupStack      i16
	sizeOfItemFlagsStack  i16
	sizeOfBeginPopupStack i16
	sizeOfDisabledStack   i16
}

struct WindowStackData {
	window                              &Window
	parentLastItemDataBackup            LastItemData
	stackSizesInBegin                   ErrorRecoveryState
	disabledOverrideReenable            bool
	disabledOverrideReenableAlphaBackup f32
}

struct ShrinkWidthItem {
	index        int
	width        f32
	initialWidth f32
}

struct PtrOrIndex {
	ptr   voidptr
	index int
}

struct DeactivatedItemData {
	iD                  ID
	elapseFrame         int
	hasBeenEditedBefore bool
	isAlive             bool
}

enum PopupPositionPolicy {
	default
	combo_box
	tooltip
}

struct PopupData {
	popupId          ID
	window           &Window
	restoreNavWindow &Window
	parentNavLayer   int
	openFrameCount   int
	openParentId     ID
	openPopupPos     ImVec2
	openMousePos     ImVec2
}

struct ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN {
	storage [5]ImU32
}

type ImBitArrayForNamedKeys = ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN

enum ImGuiInputEventType {
	none = 0
	mouse_pos
	mouse_wheel
	mouse_button
	mouse_viewport
	key
	text
	focus
	count
}

enum InputSource {
	none = 0
	mouse
	keyboard
	gamepad
	count
}

struct ImGuiInputEventMousePos {
	posX        f32
	posY        f32
	mouseSource MouseSource
}

struct ImGuiInputEventMouseWheel {
	wheelX      f32
	wheelY      f32
	mouseSource MouseSource
}

struct ImGuiInputEventMouseButton {
	button      int
	down        bool
	mouseSource MouseSource
}

struct ImGuiInputEventMouseViewport {
	hoveredViewportID ID
}

struct ImGuiInputEventKey {
	key         Key
	down        bool
	analogValue f32
}

struct ImGuiInputEventText {
	char u32
}

struct ImGuiInputEventAppFocused {
	focused bool
}

struct KeyRoutingIndex {
	type              ImGuiInputEventType
	source            InputSource
	eventId           ImU32
	addedByTestEngine bool
}

struct KeyRoutingData {
	nextEntryIndex   KeyRoutingIndex
	mods             ImU16
	routingCurrScore ImU8
	routingNextScore ImU8
	routingCurr      ID
	routingNext      ID
}

struct ImVector_ImGuiKeyRoutingData {
	size     int
	capacity int
	data     &KeyRoutingData
}

struct KeyRoutingTable {
	index       [155]KeyRoutingIndex
	entries     ImVector_ImGuiKeyRoutingData
	entriesNext ImVector_ImGuiKeyRoutingData
}

struct KeyOwnerData {
	ownerCurr        ID
	ownerNext        ID
	lockThisFrame    bool
	lockUntilRelease bool
}

enum InputFlagsPrivate_ {
	repeat_rate_default                    = 1 << 1
	repeat_rate_nav_move                   = 1 << 2
	repeat_rate_nav_tweak                  = 1 << 3
	repeat_until_release                   = 1 << 4
	repeat_until_key_mods_change           = 1 << 5
	repeat_until_key_mods_change_from_none = 1 << 6
	repeat_until_other_key_press           = 1 << 7
	lock_this_frame                        = 1 << 20
	lock_until_release                     = 1 << 21
	cond_hovered                           = 1 << 22
	cond_active                            = 1 << 23
	cond_default_                          = 1 << 22 | 1 << 23
	repeat_rate_mask_                      = 1 << 1 | 1 << 2 | 1 << 3
	repeat_until_mask_                     = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	repeat_mask_                           = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	cond_mask_                             = 1 << 22 | 1 << 23
	route_type_mask_                       = 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13
	route_options_mask_                    = 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
	supported_by_is_key_pressed            = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	supported_by_is_mouse_clicked          = 1 << 0
	supported_by_shortcut                  = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
	supported_by_set_next_item_shortcut    = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17 | 1 << 18
	supported_by_set_key_owner             = 1 << 20 | 1 << 21
	supported_by_set_item_key_owner        = 1 << 20 | 1 << 21 | 1 << 22 | 1 << 23
}

struct ListClipperRange {
	min                 int
	max                 int
	posToIndexConvert   bool
	posToIndexOffsetMin ImS8
	posToIndexOffsetMax ImS8
}

struct ImVector_ImGuiListClipperRange {
	size     int
	capacity int
	data     &ListClipperRange
}

struct ListClipperData {
	listClipper     &ListClipper
	lossynessOffset f32
	stepNo          int
	itemsFrozen     int
	ranges          ImVector_ImGuiListClipperRange
}

enum ActivateFlags_ {
	none                  = 0
	prefer_input          = 1 << 0
	prefer_tweak          = 1 << 1
	try_to_preserve_state = 1 << 2
	from_tabbing          = 1 << 3
	from_shortcut         = 1 << 4
}

enum ScrollFlags_ {
	none                  = 0
	keep_visible_edge_x   = 1 << 0
	keep_visible_edge_y   = 1 << 1
	keep_visible_center_x = 1 << 2
	keep_visible_center_y = 1 << 3
	always_center_x       = 1 << 4
	always_center_y       = 1 << 5
	no_scroll_parent      = 1 << 6
	mask_x_               = 1 << 0 | 1 << 2 | 1 << 4
	mask_y_               = 1 << 1 | 1 << 3 | 1 << 5
}

enum NavRenderCursorFlags_ {
	none        = 0
	compact     = 1 << 1
	always_draw = 1 << 2
	no_rounding = 1 << 3
}

enum NavMoveFlags_ {
	none                      = 0
	loop_x                    = 1 << 0
	loop_y                    = 1 << 1
	wrap_x                    = 1 << 2
	wrap_y                    = 1 << 3
	wrap_mask_                = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
	allow_current_nav_id      = 1 << 4
	also_score_visible_set    = 1 << 5
	scroll_to_edge_y          = 1 << 6
	forwarded                 = 1 << 7
	debug_no_result           = 1 << 8
	focus_api                 = 1 << 9
	is_tabbing                = 1 << 10
	is_page_move              = 1 << 11
	activate                  = 1 << 12
	no_select                 = 1 << 13
	no_set_nav_cursor_visible = 1 << 14
	no_clear_active_id        = 1 << 15
}

enum NavLayer {
	main = 0
	menu = 1
	count
}

struct NavItemData {
	window            &Window
	iD                ID
	focusScopeId      ID
	rectRel           C.ImRect
	itemFlags         ItemFlags
	distBox           f32
	distCenter        f32
	distAxial         f32
	selectionUserData SelectionUserData
}

struct FocusScopeData {
	iD       ID
	windowID ID
}

enum TypingSelectFlags_ {
	none                   = 0
	allow_backspace        = 1 << 0
	allow_single_char_mode = 1 << 1
}

struct TypingSelectRequest {
	flags           TypingSelectFlags
	searchBufferLen int
	searchBuffer    &i8
	selectRequest   bool
	singleCharMode  bool
	singleCharSize  ImS8
}

struct TypingSelectState {
	request            TypingSelectRequest
	searchBuffer       [64]i8
	focusScope         ID
	lastRequestFrame   int
	lastRequestTime    f32
	singleCharModeLock bool
}

enum OldColumnFlags_ {
	none                      = 0
	no_border                 = 1 << 0
	no_resize                 = 1 << 1
	no_preserve_widths        = 1 << 2
	no_force_within_window    = 1 << 3
	grow_parent_contents_size = 1 << 4
}

struct OldColumnData {
	offsetNorm             f32
	offsetNormBeforeResize f32
	flags                  OldColumnFlags
	clipRect               C.ImRect
}

struct ImVector_ImGuiOldColumnData {
	size     int
	capacity int
	data     &OldColumnData
}

struct OldColumns {
	iD                       ID
	flags                    OldColumnFlags
	isFirstFrame             bool
	isBeingResized           bool
	current                  int
	count                    int
	offMinX                  f32
	offMaxX                  f32
	lineMinY                 f32
	lineMaxY                 f32
	hostCursorPosY           f32
	hostCursorMaxPosX        f32
	hostInitialClipRect      C.ImRect
	hostBackupClipRect       C.ImRect
	hostBackupParentWorkRect C.ImRect
	columns                  ImVector_ImGuiOldColumnData
	splitter                 ImDrawListSplitter
}

struct BoxSelectState {
	iD                    ID
	isActive              bool
	isStarting            bool
	isStartedFromVoid     bool
	isStartedSetNavIdOnce bool
	requestClear          bool
	keyMods               KeyChord
	startPosRel           ImVec2
	endPosRel             ImVec2
	scrollAccum           ImVec2
	window                &Window
	unclipMode            bool
	unclipRect            C.ImRect
	boxSelectRectPrev     C.ImRect
	boxSelectRectCurr     C.ImRect
}

struct MultiSelectTempData {
	iO                 MultiSelectIO
	storage            &MultiSelectState
	focusScopeId       ID
	flags              MultiSelectFlags
	scopeRectMin       ImVec2
	backupCursorMaxPos ImVec2
	lastSubmittedItem  SelectionUserData
	boxSelectId        ID
	keyMods            KeyChord
	loopRequestSetAll  ImS8
	isEndIO            bool
	isFocused          bool
	isKeyboardSetRange bool
	navIdPassedBy      bool
	rangeSrcPassedBy   bool
	rangeDstPassedBy   bool
}

struct MultiSelectState {
	window            &Window
	iD                ID
	lastFrameActive   int
	lastSelectionSize int
	rangeSelected     ImS8
	navIdSelected     ImS8
	rangeSrcItem      SelectionUserData
	navIdItem         SelectionUserData
}

enum DockNodeFlagsPrivate_ {
	dock_space                    = 1 << 10
	central_node                  = 1 << 11
	no_tab_bar                    = 1 << 12
	hidden_tab_bar                = 1 << 13
	no_window_menu_button         = 1 << 14
	no_close_button               = 1 << 15
	no_resize_x                   = 1 << 16
	no_resize_y                   = 1 << 17
	docked_windows_in_focus_route = 1 << 18
	no_docking_split_other        = 1 << 19
	no_docking_over_me            = 1 << 20
	no_docking_over_other         = 1 << 21
	no_docking_over_empty         = 1 << 22
	no_docking                    = 1 << 20 | 1 << 21 | 1 << 22 | 1 << 4 | 1 << 19
	shared_flags_inherit_mask_    = int(~0)
	no_resize_flags_mask_         = 1 << 5 | 1 << 16 | 1 << 17
	local_flags_transfer_mask_    = 1 << 4 | 1 << 5 | 1 << 16 | 1 << 17 | 1 << 6 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15
	saved_flags_mask_             = 1 << 5 | 1 << 16 | 1 << 17 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15
}

enum DataAuthority_ {
	auto
	dock_node
	window
}

enum DockNodeState {
	unknown
	host_window_hidden_because_single_window
	host_window_hidden_because_windows_are_resizing
	host_window_visible
}

struct ImVector_ImGuiWindowPtr {
	size     int
	capacity int
	data     &&Window
}

struct DockNode {
	iD                     ID
	sharedFlags            DockNodeFlags
	localFlags             DockNodeFlags
	localFlagsInWindows    DockNodeFlags
	mergedFlags            DockNodeFlags
	state                  DockNodeState
	parentNode             &DockNode
	childNodes             [2]&DockNode
	windows                ImVector_ImGuiWindowPtr
	tabBar                 &C.ImGuiTabBar
	pos                    ImVec2
	size                   ImVec2
	sizeRef                ImVec2
	splitAxis              Axis
	windowClass            WindowClass
	lastBgColor            ImU32
	hostWindow             &Window
	visibleWindow          &Window
	centralNode            &DockNode
	onlyNodeWithWindows    &DockNode
	countNodeWithWindows   int
	lastFrameAlive         int
	lastFrameActive        int
	lastFrameFocused       int
	lastFocusedNodeId      ID
	selectedTabId          ID
	wantCloseTabId         ID
	refViewportId          ID
	authorityForPos        DataAuthority
	authorityForSize       DataAuthority
	authorityForViewport   DataAuthority
	isVisible              bool
	isFocused              bool
	isBgDrawnThisFrame     bool
	hasCloseButton         bool
	hasWindowMenuButton    bool
	hasCentralNodeChild    bool
	wantCloseAll           bool
	wantLockSizeOnce       bool
	wantMouseMove          bool
	wantHiddenTabBarUpdate bool
	wantHiddenTabBarToggle bool
}

enum WindowDockStyleCol {
	text
	tab_hovered
	tab_focused
	tab_selected
	tab_selected_overline
	tab_dimmed
	tab_dimmed_selected
	tab_dimmed_selected_overline
	count
}

struct WindowDockStyle {
	colors [8]ImU32
}

struct ImVector_ImGuiDockRequest {
	size     int
	capacity int
	data     &C.ImGuiDockRequest
}

struct ImVector_ImGuiDockNodeSettings {
	size     int
	capacity int
	data     &C.ImGuiDockNodeSettings
}

struct DockContext {
	nodes           Storage
	requests        ImVector_ImGuiDockRequest
	nodesSettings   ImVector_ImGuiDockNodeSettings
	wantFullRebuild bool
}

struct ViewportP {
	_ImGuiViewport          Viewport
	window                  &Window
	idx                     int
	lastFrameActive         int
	lastFocusedStampCount   int
	lastNameHash            ID
	lastPos                 ImVec2
	lastSize                ImVec2
	alpha                   f32
	lastAlpha               f32
	lastFocusedHadNavWindow bool
	platformMonitor         i16
	bgFgDrawListsLastFrame  [2]int
	bgFgDrawLists           [2]&ImDrawList
	drawDataP               ImDrawData
	drawDataBuilder         ImDrawDataBuilder
	lastPlatformPos         ImVec2
	lastPlatformSize        ImVec2
	lastRendererSize        ImVec2
	workInsetMin            ImVec2
	workInsetMax            ImVec2
	buildWorkInsetMin       ImVec2
	buildWorkInsetMax       ImVec2
}

struct WindowSettings {
	iD          ID
	pos         ImVec2ih
	size        ImVec2ih
	viewportPos ImVec2ih
	viewportId  ID
	dockId      ID
	classId     ID
	dockOrder   i16
	collapsed   bool
	isChild     bool
	wantApply   bool
	wantDelete  bool
}

struct SettingsHandler {
	typeName   &i8
	typeHash   ID
	clearAllFn fn (&Context, &SettingsHandler)
	readInitFn fn (&Context, &SettingsHandler)
	readOpenFn fn (&Context, &SettingsHandler, &i8) voidptr
	readLineFn fn (&Context, &SettingsHandler, voidptr, &i8)
	applyAllFn fn (&Context, &SettingsHandler)
	writeAllFn fn (&Context, &SettingsHandler, &TextBuffer)
	userData   voidptr
}

enum LocKey {
	version_str                         = 0
	table_size_one                      = 1
	table_size_all_fit                  = 2
	table_size_all_default              = 3
	table_reset_order                   = 4
	windowing_main_menu_bar             = 5
	windowing_popup                     = 6
	windowing_untitled                  = 7
	open_link_s                         = 8
	copy_link                           = 9
	docking_hide_tab_bar                = 10
	docking_hold_shift_to_dock          = 11
	docking_drag_to_undock_or_move_node = 12
	count                               = 13
}

struct ErrorCallback {
	key  LocKey
	text &i8
}

enum DebugLogFlags_ {
	none                  = 0
	event_error           = 1 << 0
	event_active_id       = 1 << 1
	event_focus           = 1 << 2
	event_popup           = 1 << 3
	event_nav             = 1 << 4
	event_clipper         = 1 << 5
	event_selection       = 1 << 6
	event_io              = 1 << 7
	event_font            = 1 << 8
	event_input_routing   = 1 << 9
	event_docking         = 1 << 10
	event_viewport        = 1 << 11
	event_mask_           = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8 | 1 << 9 | 1 << 10 | 1 << 11
	output_to_tty         = 1 << 20
	output_to_test_engine = 1 << 21
}

struct DebugAllocEntry {
	frameCount int
	allocCount ImS16
	freeCount  ImS16
}

struct DebugAllocInfo {
	totalAllocCount int
	totalFreeCount  int
	lastEntriesIdx  ImS16
	lastEntriesBuf  [6]DebugAllocEntry
}

struct MetricsConfig {
	showDebugLog             bool
	showIDStackTool          bool
	showWindowsRects         bool
	showWindowsBeginOrder    bool
	showTablesRects          bool
	showDrawCmdMesh          bool
	showDrawCmdBoundingBoxes bool
	showTextEncodingViewer   bool
	showDockingNodes         bool
	showWindowsRectsType     int
	showTablesRectsType      int
	highlightMonitorIdx      int
	highlightViewportID      ID
}

struct StackLevelInfo {
	iD              ID
	queryFrameCount ImS8
	querySuccess    bool
	dataType        DataType
	desc            [57]i8
}

struct ImVector_ImGuiStackLevelInfo {
	size     int
	capacity int
	data     &StackLevelInfo
}

struct ContextHookCallback {
	lastActiveFrame         int
	stackLevel              int
	queryId                 ID
	results                 ImVector_ImGuiStackLevelInfo
	copyToClipboardOnCtrlC  bool
	copyToClipboardLastTime f32
	resultPathBuf           TextBuffer
}

enum ContextHookType {
	new_frame_pre
	new_frame_post
	end_frame_pre
	end_frame_post
	render_pre
	render_post
	shutdown
	pending_removal_
}

struct ContextHook {
	hookId   ID
	type     ContextHookType
	owner    ID
	callback ContextHookCallback
	userData voidptr
}

struct ImVector_ImGuiInputEvent {
	size     int
	capacity int
	data     &C.ImGuiInputEvent
}

struct ImVector_ImGuiWindowStackData {
	size     int
	capacity int
	data     &WindowStackData
}

struct ImVector_ImGuiColorMod {
	size     int
	capacity int
	data     &ColorMod
}

struct ImVector_ImGuiStyleMod {
	size     int
	capacity int
	data     &StyleMod
}

struct ImVector_ImGuiFocusScopeData {
	size     int
	capacity int
	data     &FocusScopeData
}

struct ImVector_ImGuiItemFlags {
	size     int
	capacity int
	data     &ItemFlags
}

struct ImVector_ImGuiGroupData {
	size     int
	capacity int
	data     &GroupData
}

struct ImVector_ImGuiPopupData {
	size     int
	capacity int
	data     &PopupData
}

struct ImVector_ImGuiTreeNodeStackData {
	size     int
	capacity int
	data     &TreeNodeStackData
}

struct ImVector_ImGuiViewportPPtr {
	size     int
	capacity int
	data     &&ViewportP
}

struct ImVector_unsigned_char {
	size     int
	capacity int
	data     &u8
}

struct ImVector_ImGuiListClipperData {
	size     int
	capacity int
	data     &ListClipperData
}

struct ImVector_ImGuiTableTempData {
	size     int
	capacity int
	data     &TableTempData
}

struct ImVector_ImGuiTable {
	size     int
	capacity int
	data     &Table
}

struct ImPool_ImGuiTable {
	buf        ImVector_ImGuiTable
	map        Storage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImGuiTabBar {
	size     int
	capacity int
	data     &C.ImGuiTabBar
}

struct ImPool_ImGuiTabBar {
	buf        ImVector_ImGuiTabBar
	map        Storage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImGuiPtrOrIndex {
	size     int
	capacity int
	data     &PtrOrIndex
}

struct ImVector_ImGuiShrinkWidthItem {
	size     int
	capacity int
	data     &ShrinkWidthItem
}

struct ImVector_ImGuiMultiSelectTempData {
	size     int
	capacity int
	data     &MultiSelectTempData
}

struct ImVector_ImGuiMultiSelectState {
	size     int
	capacity int
	data     &MultiSelectState
}

struct ImPool_ImGuiMultiSelectState {
	buf        ImVector_ImGuiMultiSelectState
	map        Storage
	freeIdx    ImPoolIdx
	aliveCount ImPoolIdx
}

struct ImVector_ImGuiID {
	size     int
	capacity int
	data     &ID
}

struct ImVector_ImGuiSettingsHandler {
	size     int
	capacity int
	data     &SettingsHandler
}

struct ImChunkStream_ImGuiWindowSettings {
	buf ImVector_char
}

struct ImChunkStream_ImGuiTableSettings {
	buf ImVector_char
}

struct ImVector_ImGuiContextHook {
	size     int
	capacity int
	data     &ContextHook
}

struct Context {
	initialized                        bool
	fontAtlasOwnedByContext            bool
	iO                                 IO
	platformIO                         PlatformIO
	style                              Style
	configFlagsCurrFrame               ConfigFlags
	configFlagsLastFrame               ConfigFlags
	font                               &ImFont
	fontSize                           f32
	fontBaseSize                       f32
	fontScale                          f32
	currentDpiScale                    f32
	drawListSharedData                 ImDrawListSharedData
	time                               f64
	frameCount                         int
	frameCountEnded                    int
	frameCountPlatformEnded            int
	frameCountRendered                 int
	withinEndChildID                   ID
	withinFrameScope                   bool
	withinFrameScopeWithImplicitWindow bool
	gcCompactAll                       bool
	testEngineHookItems                bool
	testEngine                         voidptr
	contextName                        [16]i8
	inputEventsQueue                   ImVector_ImGuiInputEvent
	inputEventsTrail                   ImVector_ImGuiInputEvent
	inputEventsNextMouseSource         MouseSource
	inputEventsNextEventId             ImU32
	windows                            ImVector_ImGuiWindowPtr
	windowsFocusOrder                  ImVector_ImGuiWindowPtr
	windowsTempSortBuffer              ImVector_ImGuiWindowPtr
	currentWindowStack                 ImVector_ImGuiWindowStackData
	windowsById                        Storage
	windowsActiveCount                 int
	windowsBorderHoverPadding          f32
	debugBreakInWindow                 ID
	currentWindow                      &Window
	hoveredWindow                      &Window
	hoveredWindowUnderMovingWindow     &Window
	hoveredWindowBeforeClear           &Window
	movingWindow                       &Window
	wheelingWindow                     &Window
	wheelingWindowRefMousePos          ImVec2
	wheelingWindowStartFrame           int
	wheelingWindowScrolledFrame        int
	wheelingWindowReleaseTimer         f32
	wheelingWindowWheelRemainder       ImVec2
	wheelingAxisAvg                    ImVec2
	debugDrawIdConflicts               ID
	debugHookIdInfo                    ID
	hoveredId                          ID
	hoveredIdPreviousFrame             ID
	hoveredIdPreviousFrameItemCount    int
	hoveredIdTimer                     f32
	hoveredIdNotActiveTimer            f32
	hoveredIdAllowOverlap              bool
	hoveredIdIsDisabled                bool
	itemUnclipByLog                    bool
	activeId                           ID
	activeIdIsAlive                    ID
	activeIdTimer                      f32
	activeIdIsJustActivated            bool
	activeIdAllowOverlap               bool
	activeIdNoClearOnFocusLoss         bool
	activeIdHasBeenPressedBefore       bool
	activeIdHasBeenEditedBefore        bool
	activeIdHasBeenEditedThisFrame     bool
	activeIdFromShortcut               bool
	activeIdMouseButton                int
	activeIdClickOffset                ImVec2
	activeIdWindow                     &Window
	activeIdSource                     InputSource
	activeIdPreviousFrame              ID
	deactivatedItemData                DeactivatedItemData
	activeIdValueOnActivation          DataTypeStorage
	lastActiveId                       ID
	lastActiveIdTimer                  f32
	lastKeyModsChangeTime              f64
	lastKeyModsChangeFromNoneTime      f64
	lastKeyboardKeyPressTime           f64
	keysMayBeCharInput                 ImBitArrayForNamedKeys
	keysOwnerData                      [155]KeyOwnerData
	keysRoutingTable                   KeyRoutingTable
	activeIdUsingNavDirMask            ImU32
	activeIdUsingAllKeyboardKeys       bool
	debugBreakInShortcutRouting        KeyChord
	currentFocusScopeId                ID
	currentItemFlags                   ItemFlags
	debugLocateId                      ID
	nextItemData                       NextItemData
	lastItemData                       LastItemData
	nextWindowData                     NextWindowData
	debugShowGroupRects                bool
	debugFlashStyleColorIdx            Col
	colorStack                         ImVector_ImGuiColorMod
	styleVarStack                      ImVector_ImGuiStyleMod
	fontStack                          ImVector_ImFontPtr
	focusScopeStack                    ImVector_ImGuiFocusScopeData
	itemFlagsStack                     ImVector_ImGuiItemFlags
	groupStack                         ImVector_ImGuiGroupData
	openPopupStack                     ImVector_ImGuiPopupData
	beginPopupStack                    ImVector_ImGuiPopupData
	treeNodeStack                      ImVector_ImGuiTreeNodeStackData
	viewports                          ImVector_ImGuiViewportPPtr
	currentViewport                    &ViewportP
	mouseViewport                      &ViewportP
	mouseLastHoveredViewport           &ViewportP
	platformLastFocusedViewportId      ID
	fallbackMonitor                    PlatformMonitor
	platformMonitorsFullWorkRect       C.ImRect
	viewportCreatedCount               int
	platformWindowsCreatedCount        int
	viewportFocusedStampCount          int
	navCursorVisible                   bool
	navHighlightItemUnderNav           bool
	navMousePosDirty                   bool
	navIdIsAlive                       bool
	navId                              ID
	navWindow                          &Window
	navFocusScopeId                    ID
	navLayer                           NavLayer
	navActivateId                      ID
	navActivateDownId                  ID
	navActivatePressedId               ID
	navActivateFlags                   ActivateFlags
	navFocusRoute                      ImVector_ImGuiFocusScopeData
	navHighlightActivatedId            ID
	navHighlightActivatedTimer         f32
	navNextActivateId                  ID
	navNextActivateFlags               ActivateFlags
	navInputSource                     InputSource
	navLastValidSelectionUserData      SelectionUserData
	navCursorHideFrames                ImS8
	navAnyRequest                      bool
	navInitRequest                     bool
	navInitRequestFromMove             bool
	navInitResult                      NavItemData
	navMoveSubmitted                   bool
	navMoveScoringItems                bool
	navMoveForwardToNextFrame          bool
	navMoveFlags                       NavMoveFlags
	navMoveScrollFlags                 ScrollFlags
	navMoveKeyMods                     KeyChord
	navMoveDir                         Dir
	navMoveDirForDebug                 Dir
	navMoveClipDir                     Dir
	navScoringRect                     C.ImRect
	navScoringNoClipRect               C.ImRect
	navScoringDebugCount               int
	navTabbingDir                      int
	navTabbingCounter                  int
	navMoveResultLocal                 NavItemData
	navMoveResultLocalVisible          NavItemData
	navMoveResultOther                 NavItemData
	navTabbingResultFirst              NavItemData
	navJustMovedFromFocusScopeId       ID
	navJustMovedToId                   ID
	navJustMovedToFocusScopeId         ID
	navJustMovedToKeyMods              KeyChord
	navJustMovedToIsTabbing            bool
	navJustMovedToHasSelectionData     bool
	configNavWindowingKeyNext          KeyChord
	configNavWindowingKeyPrev          KeyChord
	navWindowingTarget                 &Window
	navWindowingTargetAnim             &Window
	navWindowingListWindow             &Window
	navWindowingTimer                  f32
	navWindowingHighlightAlpha         f32
	navWindowingToggleLayer            bool
	navWindowingToggleKey              Key
	navWindowingAccumDeltaPos          ImVec2
	navWindowingAccumDeltaSize         ImVec2
	dimBgRatio                         f32
	dragDropActive                     bool
	dragDropWithinSource               bool
	dragDropWithinTarget               bool
	dragDropSourceFlags                DragDropFlags
	dragDropSourceFrameCount           int
	dragDropMouseButton                int
	dragDropPayload                    Payload
	dragDropTargetRect                 C.ImRect
	dragDropTargetClipRect             C.ImRect
	dragDropTargetId                   ID
	dragDropAcceptFlags                DragDropFlags
	dragDropAcceptIdCurrRectSurface    f32
	dragDropAcceptIdCurr               ID
	dragDropAcceptIdPrev               ID
	dragDropAcceptFrameCount           int
	dragDropHoldJustPressedId          ID
	dragDropPayloadBufHeap             ImVector_unsigned_char
	dragDropPayloadBufLocal            [16]u8
	clipperTempDataStacked             int
	clipperTempData                    ImVector_ImGuiListClipperData
	currentTable                       &Table
	debugBreakInTable                  ID
	tablesTempDataStacked              int
	tablesTempData                     ImVector_ImGuiTableTempData
	tables                             ImPool_ImGuiTable
	tablesLastTimeActive               ImVector_float
	drawChannelsTempMergeBuffer        ImVector_ImDrawChannel
	currentTabBar                      &C.ImGuiTabBar
	tabBars                            ImPool_ImGuiTabBar
	currentTabBarStack                 ImVector_ImGuiPtrOrIndex
	shrinkWidthBuffer                  ImVector_ImGuiShrinkWidthItem
	boxSelectState                     BoxSelectState
	currentMultiSelect                 &MultiSelectTempData
	multiSelectTempDataStacked         int
	multiSelectTempData                ImVector_ImGuiMultiSelectTempData
	multiSelectStorage                 ImPool_ImGuiMultiSelectState
	hoverItemDelayId                   ID
	hoverItemDelayIdPreviousFrame      ID
	hoverItemDelayTimer                f32
	hoverItemDelayClearTimer           f32
	hoverItemUnlockedStationaryId      ID
	hoverWindowUnlockedStationaryId    ID
	mouseCursor                        MouseCursor
	mouseStationaryTimer               f32
	mouseLastValidPos                  ImVec2
	inputTextState                     InputTextState
	inputTextDeactivatedState          InputTextDeactivatedState
	inputTextPasswordFont              ImFont
	tempInputId                        ID
	dataTypeZeroValue                  DataTypeStorage
	beginMenuDepth                     int
	beginComboDepth                    int
	colorEditOptions                   ColorEditFlags
	colorEditCurrentID                 ID
	colorEditSavedID                   ID
	colorEditSavedHue                  f32
	colorEditSavedSat                  f32
	colorEditSavedColor                ImU32
	colorPickerRef                     C.ImVec4
	comboPreviewData                   ComboPreviewData
	windowResizeBorderExpectedRect     C.ImRect
	windowResizeRelativeMode           bool
	scrollbarSeekMode                  i16
	scrollbarClickDeltaToGrabCenter    f32
	sliderGrabClickOffset              f32
	sliderCurrentAccum                 f32
	sliderCurrentAccumDirty            bool
	dragCurrentAccumDirty              bool
	dragCurrentAccum                   f32
	dragSpeedDefaultRatio              f32
	disabledAlphaBackup                f32
	disabledStackSize                  i16
	tooltipOverrideCount               i16
	tooltipPreviousWindow              &Window
	clipboardHandlerData               ImVector_char
	menusIdSubmittedThisFrame          ImVector_ImGuiID
	typingSelectState                  TypingSelectState
	platformImeData                    PlatformImeData
	platformImeDataPrev                PlatformImeData
	platformImeViewport                ID
	dockContext                        DockContext
	dockNodeWindowMenuHandler          fn (&Context, &DockNode, &C.ImGuiTabBar)
	settingsLoaded                     bool
	settingsDirtyTimer                 f32
	settingsIniData                    TextBuffer
	settingsHandlers                   ImVector_ImGuiSettingsHandler
	settingsWindows                    ImChunkStream_ImGuiWindowSettings
	settingsTables                     ImChunkStream_ImGuiTableSettings
	hooks                              ImVector_ImGuiContextHook
	hookIdNext                         ID
	localizationTable                  [13]&i8
	logEnabled                         bool
	logFlags                           LogFlags
	logWindow                          &Window
	logFile                            ImFileHandle
	logBuffer                          TextBuffer
	logNextPrefix                      &i8
	logNextSuffix                      &i8
	logLinePosY                        f32
	logLineFirstItem                   bool
	logDepthRef                        int
	logDepthToExpand                   int
	logDepthToExpandDefault            int
	errorCallback                      ErrorCallback
	errorCallbackUserData              voidptr
	errorTooltipLockedPos              ImVec2
	errorFirst                         bool
	errorCountCurrentFrame             int
	stackSizesInNewFrame               ErrorRecoveryState
	stackSizesInBeginForCurrentWindow  &ErrorRecoveryState
	debugDrawIdConflictsCount          int
	debugLogFlags                      DebugLogFlags
	debugLogBuf                        TextBuffer
	debugLogIndex                      TextIndex
	debugLogSkippedErrors              int
	debugLogAutoDisableFlags           DebugLogFlags
	debugLogAutoDisableFrames          ImU8
	debugLocateFrames                  ImU8
	debugBreakInLocateId               bool
	debugBreakKeyChord                 KeyChord
	debugBeginReturnValueCullDepth     ImS8
	debugItemPickerActive              bool
	debugItemPickerMouseButton         ImU8
	debugItemPickerBreakId             ID
	debugFlashStyleColorTime           f32
	debugFlashStyleColorBackup         C.ImVec4
	debugMetricsConfig                 MetricsConfig
	debugIDStackTool                   C.ImGuiIDStackTool
	debugAllocInfo                     DebugAllocInfo
	debugHoveredDockNode               &DockNode
	framerateSecPerFrame               [60]f32
	framerateSecPerFrameIdx            int
	framerateSecPerFrameCount          int
	framerateSecPerFrameAccum          f32
	wantCaptureMouseNextFrame          int
	wantCaptureKeyboardNextFrame       int
	wantTextInputNextFrame             int
	tempBuffer                         ImVector_char
	tempKeychordName                   [64]i8
}

struct WindowTempData {
	cursorPos                 ImVec2
	cursorPosPrevLine         ImVec2
	cursorStartPos            ImVec2
	cursorMaxPos              ImVec2
	idealMaxPos               ImVec2
	currLineSize              ImVec2
	prevLineSize              ImVec2
	currLineTextBaseOffset    f32
	prevLineTextBaseOffset    f32
	isSameLine                bool
	isSetPos                  bool
	indent                    ImVec1
	columnsOffset             ImVec1
	groupOffset               ImVec1
	cursorStartPosLossyness   ImVec2
	navLayerCurrent           NavLayer
	navLayersActiveMask       i16
	navLayersActiveMaskNext   i16
	navIsScrollPushableX      bool
	navHideHighlightOneFrame  bool
	navWindowHasScrollY       bool
	menuBarAppending          bool
	menuBarOffset             ImVec2
	menuColumns               MenuColumns
	treeDepth                 int
	treeHasStackDataDepthMask ImU32
	childWindows              ImVector_ImGuiWindowPtr
	stateStorage              &Storage
	currentColumns            &OldColumns
	currentTableIdx           int
	layoutType                LayoutType
	parentLayoutType          LayoutType
	modalDimBgColor           ImU32
	windowItemStatusFlags     ItemStatusFlags
	childItemStatusFlags      ItemStatusFlags
	dockTabItemStatusFlags    ItemStatusFlags
	dockTabItemRect           C.ImRect
	itemWidth                 f32
	textWrapPos               f32
	itemWidthStack            ImVector_float
	textWrapPosStack          ImVector_float
}

struct ImVector_ImGuiOldColumns {
	size     int
	capacity int
	data     &OldColumns
}

struct Window {
	ctx                                &Context
	name                               &i8
	iD                                 ID
	flags                              WindowFlags
	flagsPreviousFrame                 WindowFlags
	childFlags                         ChildFlags
	windowClass                        WindowClass
	viewport                           &ViewportP
	viewportId                         ID
	viewportPos                        ImVec2
	viewportAllowPlatformMonitorExtend int
	pos                                ImVec2
	size                               ImVec2
	sizeFull                           ImVec2
	contentSize                        ImVec2
	contentSizeIdeal                   ImVec2
	contentSizeExplicit                ImVec2
	windowPadding                      ImVec2
	windowRounding                     f32
	windowBorderSize                   f32
	titleBarHeight                     f32
	menuBarHeight                      f32
	decoOuterSizeX1                    f32
	decoOuterSizeY1                    f32
	decoOuterSizeX2                    f32
	decoOuterSizeY2                    f32
	decoInnerSizeX1                    f32
	decoInnerSizeY1                    f32
	nameBufLen                         int
	moveId                             ID
	tabId                              ID
	childId                            ID
	popupId                            ID
	scroll                             ImVec2
	scrollMax                          ImVec2
	scrollTarget                       ImVec2
	scrollTargetCenterRatio            ImVec2
	scrollTargetEdgeSnapDist           ImVec2
	scrollbarSizes                     ImVec2
	scrollbarX                         bool
	scrollbarY                         bool
	scrollbarXStabilizeEnabled         bool
	scrollbarXStabilizeToggledHistory  ImU8
	viewportOwned                      bool
	active                             bool
	wasActive                          bool
	writeAccessed                      bool
	collapsed                          bool
	wantCollapseToggle                 bool
	skipItems                          bool
	skipRefresh                        bool
	appearing                          bool
	hidden                             bool
	isFallbackWindow                   bool
	isExplicitChild                    bool
	hasCloseButton                     bool
	resizeBorderHovered                i8
	resizeBorderHeld                   i8
	beginCount                         i16
	beginCountPreviousFrame            i16
	beginOrderWithinParent             i16
	beginOrderWithinContext            i16
	focusOrder                         i16
	autoFitFramesX                     ImS8
	autoFitFramesY                     ImS8
	autoFitOnlyGrows                   bool
	autoPosLastDirection               Dir
	hiddenFramesCanSkipItems           ImS8
	hiddenFramesCannotSkipItems        ImS8
	hiddenFramesForRenderOnly          ImS8
	disableInputsFrames                ImS8
	setWindowPosAllowFlags             Cond
	setWindowSizeAllowFlags            Cond
	setWindowCollapsedAllowFlags       Cond
	setWindowDockAllowFlags            Cond
	setWindowPosVal                    ImVec2
	setWindowPosPivot                  ImVec2
	iDStack                            ImVector_ImGuiID
	dC                                 WindowTempData
	outerRectClipped                   C.ImRect
	innerRect                          C.ImRect
	innerClipRect                      C.ImRect
	workRect                           C.ImRect
	parentWorkRect                     C.ImRect
	clipRect                           C.ImRect
	contentRegionRect                  C.ImRect
	hitTestHoleSize                    ImVec2ih
	hitTestHoleOffset                  ImVec2ih
	lastFrameActive                    int
	lastFrameJustFocused               int
	lastTimeActive                     f32
	itemWidthDefault                   f32
	stateStorage                       Storage
	columnsStorage                     ImVector_ImGuiOldColumns
	fontWindowScale                    f32
	fontWindowScaleParents             f32
	fontDpiScale                       f32
	fontRefSize                        f32
	settingsOffset                     int
	drawList                           &ImDrawList
	drawListInst                       ImDrawList
	parentWindow                       &Window
	parentWindowInBeginStack           &Window
	rootWindow                         &Window
	rootWindowPopupTree                &Window
	rootWindowDockTree                 &Window
	rootWindowForTitleBarHighlight     &Window
	rootWindowForNav                   &Window
	parentWindowForFocusRoute          &Window
	navLastChildNavWindow              &Window
	navLastIds                         [2]ID
	navRectRel                         [2]C.ImRect
	navPreferredScoringPosRel          [2]ImVec2
	navRootFocusScopeId                ID
	memoryDrawListIdxCapacity          int
	memoryDrawListVtxCapacity          int
	memoryCompacted                    bool
	dockIsActive                       bool
	dockNodeIsVisible                  bool
	dockTabIsVisible                   bool
	dockTabWantClose                   bool
	dockOrder                          i16
	dockStyle                          WindowDockStyle
	dockNode                           &DockNode
	dockNodeAsHost                     &DockNode
	dockId                             ID
}

enum ImGuiTabBarFlagsPrivate_ {
	dock_node     = 1 << 20
	is_focused    = 1 << 21
	save_settings = 1 << 22
}

enum TabItemFlagsPrivate_ {
	section_mask_   = 1 << 6 | 1 << 7
	no_close_button = 1 << 20
	button          = 1 << 21
	invisible       = 1 << 22
	unsorted        = 1 << 23
}

struct TabItem {
	iD                ID
	flags             TabItemFlags
	window            &Window
	lastFrameVisible  int
	lastFrameSelected int
	offset            f32
	width             f32
	contentWidth      f32
	requestedWidth    f32
	nameOffset        ImS32
	beginOrder        ImS16
	indexDuringLayout ImS16
	wantClose         bool
}

struct ImVector_ImGuiTabItem {
	size     int
	capacity int
	data     &TabItem
}

struct TableColumnIdx {
	window                          &Window
	tabs                            ImVector_ImGuiTabItem
	flags                           ImGuiTabBarFlags
	iD                              ID
	selectedTabId                   ID
	nextSelectedTabId               ID
	visibleTabId                    ID
	currFrameVisible                int
	prevFrameVisible                int
	barRect                         C.ImRect
	currTabsContentsHeight          f32
	prevTabsContentsHeight          f32
	widthAllTabs                    f32
	widthAllTabsIdeal               f32
	scrollingAnim                   f32
	scrollingTarget                 f32
	scrollingTargetDistToVisibility f32
	scrollingSpeed                  f32
	scrollingRectMinX               f32
	scrollingRectMaxX               f32
	separatorMinX                   f32
	separatorMaxX                   f32
	reorderRequestTabId             ID
	reorderRequestOffset            ImS16
	beginCount                      ImS8
	wantLayout                      bool
	visibleTabWasSubmitted          bool
	tabsAddedNew                    bool
	tabsActiveCount                 ImS16
	lastTabItemIdx                  ImS16
	itemSpacingY                    f32
	framePadding                    ImVec2
	backupCursorPos                 ImVec2
	tabsNames                       TextBuffer
}

type TableDrawChannelIdx = u16

struct TableColumn {
	flags                    TableColumnFlags
	widthGiven               f32
	minX                     f32
	maxX                     f32
	widthRequest             f32
	widthAuto                f32
	widthMax                 f32
	stretchWeight            f32
	initStretchWeightOrWidth f32
	clipRect                 C.ImRect
	userID                   ID
	workMinX                 f32
	workMaxX                 f32
	itemWidth                f32
	contentMaxXFrozen        f32
	contentMaxXUnfrozen      f32
	contentMaxXHeadersUsed   f32
	contentMaxXHeadersIdeal  f32
	nameOffset               ImS16
	displayOrder             TableColumnIdx
	indexWithinEnabledSet    TableColumnIdx
	prevEnabledColumn        TableColumnIdx
	nextEnabledColumn        TableColumnIdx
	sortOrder                TableColumnIdx
	drawChannelCurrent       TableDrawChannelIdx
	drawChannelFrozen        TableDrawChannelIdx
	drawChannelUnfrozen      TableDrawChannelIdx
	isEnabled                bool
	isUserEnabled            bool
	isUserEnabledNextFrame   bool
	isVisibleX               bool
	isVisibleY               bool
	isRequestOutput          bool
	isSkipItems              bool
	isPreserveWidthAuto      bool
	navLayerCurrent          ImS8
	autoFitQueue             ImU8
	cannotSkipItemsQueue     ImU8
	sortDirection            ImU8
	sortDirectionsAvailCount ImU8
	sortDirectionsAvailMask  ImU8
	sortDirectionsAvailList  ImU8
}

struct TableCellData {
	bgColor ImU32
	column  TableColumnIdx
}

struct TableHeaderData {
	index     TableColumnIdx
	textColor ImU32
	bgColor0  ImU32
	bgColor1  ImU32
}

struct TableInstanceData {
	tableInstanceID         ID
	lastOuterHeight         f32
	lastTopHeadersRowHeight f32
	lastFrozenHeight        f32
	hoveredRowLast          int
	hoveredRowNext          int
}

struct ImSpan_ImGuiTableColumn {
	data    &TableColumn
	dataEnd &TableColumn
}

struct ImSpan_ImGuiTableColumnIdx {
	data    &TableColumnIdx
	dataEnd &TableColumnIdx
}

struct ImSpan_ImGuiTableCellData {
	data    &TableCellData
	dataEnd &TableCellData
}

struct ImVector_ImGuiTableInstanceData {
	size     int
	capacity int
	data     &TableInstanceData
}

struct ImVector_ImGuiTableColumnSortSpecs {
	size     int
	capacity int
	data     &TableColumnSortSpecs
}

struct Table {
	iD                         ID
	flags                      TableFlags
	rawData                    voidptr
	tempData                   &TableTempData
	columns                    ImSpan_ImGuiTableColumn
	displayOrderToIndex        ImSpan_ImGuiTableColumnIdx
	rowCellData                ImSpan_ImGuiTableCellData
	enabledMaskByDisplayOrder  ImBitArrayPtr
	enabledMaskByIndex         ImBitArrayPtr
	visibleMaskByIndex         ImBitArrayPtr
	settingsLoadedFlags        TableFlags
	settingsOffset             int
	lastFrameActive            int
	columnsCount               int
	currentRow                 int
	currentColumn              int
	instanceCurrent            ImS16
	instanceInteracted         ImS16
	rowPosY1                   f32
	rowPosY2                   f32
	rowMinHeight               f32
	rowCellPaddingY            f32
	rowTextBaseline            f32
	rowIndentOffsetX           f32
	rowFlags                   TableRowFlags
	lastRowFlags               TableRowFlags
	rowBgColorCounter          int
	rowBgColor                 [2]ImU32
	borderColorStrong          ImU32
	borderColorLight           ImU32
	borderX1                   f32
	borderX2                   f32
	hostIndentX                f32
	minColumnWidth             f32
	outerPaddingX              f32
	cellPaddingX               f32
	cellSpacingX1              f32
	cellSpacingX2              f32
	innerWidth                 f32
	columnsGivenWidth          f32
	columnsAutoFitWidth        f32
	columnsStretchSumWeights   f32
	resizedColumnNextWidth     f32
	resizeLockMinContentsX2    f32
	refScale                   f32
	angledHeadersHeight        f32
	angledHeadersSlope         f32
	outerRect                  C.ImRect
	innerRect                  C.ImRect
	workRect                   C.ImRect
	innerClipRect              C.ImRect
	bgClipRect                 C.ImRect
	bg0ClipRectForDrawCmd      C.ImRect
	bg2ClipRectForDrawCmd      C.ImRect
	hostClipRect               C.ImRect
	hostBackupInnerClipRect    C.ImRect
	outerWindow                &Window
	innerWindow                &Window
	columnsNames               TextBuffer
	drawSplitter               &ImDrawListSplitter
	instanceDataFirst          TableInstanceData
	instanceDataExtra          ImVector_ImGuiTableInstanceData
	sortSpecsSingle            TableColumnSortSpecs
	sortSpecsMulti             ImVector_ImGuiTableColumnSortSpecs
	sortSpecs                  TableSortSpecs
	sortSpecsCount             TableColumnIdx
	columnsEnabledCount        TableColumnIdx
	columnsEnabledFixedCount   TableColumnIdx
	declColumnsCount           TableColumnIdx
	angledHeadersCount         TableColumnIdx
	hoveredColumnBody          TableColumnIdx
	hoveredColumnBorder        TableColumnIdx
	highlightColumnHeader      TableColumnIdx
	autoFitSingleColumn        TableColumnIdx
	resizedColumn              TableColumnIdx
	lastResizedColumn          TableColumnIdx
	heldHeaderColumn           TableColumnIdx
	reorderColumn              TableColumnIdx
	reorderColumnDir           TableColumnIdx
	leftMostEnabledColumn      TableColumnIdx
	rightMostEnabledColumn     TableColumnIdx
	leftMostStretchedColumn    TableColumnIdx
	rightMostStretchedColumn   TableColumnIdx
	contextPopupColumn         TableColumnIdx
	freezeRowsRequest          TableColumnIdx
	freezeRowsCount            TableColumnIdx
	freezeColumnsRequest       TableColumnIdx
	freezeColumnsCount         TableColumnIdx
	rowCellDataCurrent         TableColumnIdx
	dummyDrawChannel           TableDrawChannelIdx
	bg2DrawChannelCurrent      TableDrawChannelIdx
	bg2DrawChannelUnfrozen     TableDrawChannelIdx
	navLayer                   ImS8
	isLayoutLocked             bool
	isInsideRow                bool
	isInitializing             bool
	isSortSpecsDirty           bool
	isUsingHeaders             bool
	isContextPopupOpen         bool
	disableDefaultContextMenu  bool
	isSettingsRequestLoad      bool
	isSettingsDirty            bool
	isDefaultDisplayOrder      bool
	isResetAllRequest          bool
	isResetDisplayOrderRequest bool
	isUnfrozenRows             bool
	isDefaultSizingPolicy      bool
	isActiveIdAliveBeforeTable bool
	isActiveIdInTable          bool
	hasScrollbarYCurr          bool
	hasScrollbarYPrev          bool
	memoryCompacted            bool
	hostSkipItems              bool
}

struct ImVector_ImGuiTableHeaderData {
	size     int
	capacity int
	data     &TableHeaderData
}

struct TableTempData {
	tableIndex                   int
	lastTimeActive               f32
	angledHeadersExtraWidth      f32
	angledHeadersRequests        ImVector_ImGuiTableHeaderData
	userOuterSize                ImVec2
	drawSplitter                 ImDrawListSplitter
	hostBackupWorkRect           C.ImRect
	hostBackupParentWorkRect     C.ImRect
	hostBackupPrevLineSize       ImVec2
	hostBackupCurrLineSize       ImVec2
	hostBackupCursorMaxPos       ImVec2
	hostBackupColumnsOffset      ImVec1
	hostBackupItemWidth          f32
	hostBackupItemWidthStackSize int
}

struct TableColumnSettings {
	widthOrWeight f32
	userID        ID
	index         TableColumnIdx
	displayOrder  TableColumnIdx
	sortOrder     TableColumnIdx
	sortDirection ImU8
	isEnabled     ImS8
	isStretch     ImU8
}

struct TableSettings {
	iD              ID
	saveFlags       TableFlags
	refScale        f32
	columnsCount    TableColumnIdx
	columnsCountMax TableColumnIdx
	wantApply       bool
}

struct ImFontBuilderIO {
	fontBuilder_Build fn (&ImFontAtlas) bool
}

// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
@[c: 'ImVec2_ImVec2_Nil']
fn im_vec2_im_vec2_nil() &ImVec2

@[c: 'ImVec2_ImVec2_Nil_Construct']
fn im_vec2_im_vec2_nil_construct(self &ImVec2)

@[c: 'ImVec2_destroy']
fn im_vec2_destroy(self &ImVec2)

@[c: 'ImVec2_ImVec2_Float']
fn im_vec2_im_vec2_float(_x f32, _y f32) &ImVec2

@[c: 'ImVec2_ImVec2_Float_Construct']
fn im_vec2_im_vec2_float_construct(self &ImVec2, _x f32, _y f32)

@[c: 'ImVec4_ImVec4_Nil']
fn im_vec4_im_vec4_nil() &C.ImVec4

@[c: 'ImVec4_ImVec4_Nil_Construct']
fn im_vec4_im_vec4_nil_construct(self &C.ImVec4)

@[c: 'ImVec4_destroy']
fn im_vec4_destroy(self &C.ImVec4)

@[c: 'ImVec4_ImVec4_Float']
fn im_vec4_im_vec4_float(_x f32, _y f32, _z f32, _w f32) &C.ImVec4

@[c: 'ImVec4_ImVec4_Float_Construct']
fn im_vec4_im_vec4_float_construct(self &C.ImVec4, _x f32, _y f32, _z f32, _w f32)

@[c: 'igCreateContext']
fn create_context(shared_font_atlas &ImFontAtlas) &Context

@[c: 'igDestroyContext']
fn destroy_context(ctx &Context)

@[c: 'igGetCurrentContext']
fn get_current_context() &Context

@[c: 'igSetCurrentContext']
fn set_current_context(ctx &Context)

@[c: 'igGetIO_Nil']
fn get_io_nil() &IO

@[c: 'igGetPlatformIO_Nil']
fn get_platform_io_nil() &PlatformIO

@[c: 'igGetStyle']
fn get_style() &Style

@[c: 'igNewFrame']
fn new_frame()

@[c: 'igEndFrame']
fn end_frame()

@[c: 'igRender']
fn render()

@[c: 'igGetDrawData']
fn get_draw_data() &ImDrawData

@[c: 'igShowDemoWindow']
fn show_demo_window(p_open &bool)

@[c: 'igShowMetricsWindow']
fn show_metrics_window(p_open &bool)

@[c: 'igShowDebugLogWindow']
fn show_debug_log_window(p_open &bool)

@[c: 'igShowIDStackToolWindow']
fn show_ids_tack_tool_window(p_open &bool)

@[c: 'igShowAboutWindow']
fn show_about_window(p_open &bool)

@[c: 'igShowStyleEditor']
fn show_style_editor(ref &Style)

@[c: 'igShowStyleSelector']
fn show_style_selector(label &i8) bool

@[c: 'igShowFontSelector']
fn show_font_selector(label &i8)

@[c: 'igShowUserGuide']
fn show_user_guide()

@[c: 'igGetVersion']
fn get_version() &i8

@[c: 'igStyleColorsDark']
fn style_colors_dark(dst &Style)

@[c: 'igStyleColorsLight']
fn style_colors_light(dst &Style)

@[c: 'igStyleColorsClassic']
fn style_colors_classic(dst &Style)

@[c: 'igBegin']
fn begin(name &i8, p_open &bool, flags WindowFlags) bool

@[c: 'igEnd']
fn end()

@[c: 'igBeginChild_Str']
fn begin_child_str(str_id &i8, size ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c: 'igBeginChild_ID']
fn begin_child_id(id ID, size ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c: 'igEndChild']
fn end_child()

@[c: 'igIsWindowAppearing']
fn is_window_appearing() bool

@[c: 'igIsWindowCollapsed']
fn is_window_collapsed() bool

@[c: 'igIsWindowFocused']
fn is_window_focused(flags FocusedFlags) bool

@[c: 'igIsWindowHovered']
fn is_window_hovered(flags HoveredFlags) bool

@[c: 'igGetWindowDrawList']
fn get_window_draw_list() &ImDrawList

@[c: 'igGetWindowDpiScale']
fn get_window_dpi_scale() f32

@[c: 'igGetWindowPos']
fn get_window_pos(p_out &ImVec2)

@[c: 'igGetWindowSize']
fn get_window_size(p_out &ImVec2)

@[c: 'igGetWindowWidth']
fn get_window_width() f32

@[c: 'igGetWindowHeight']
fn get_window_height() f32

@[c: 'igGetWindowViewport']
fn get_window_viewport() &Viewport

@[c: 'igSetNextWindowPos']
fn set_next_window_pos(pos ImVec2, cond Cond, pivot ImVec2)

@[c: 'igSetNextWindowSize']
fn set_next_window_size(size ImVec2, cond Cond)

@[c: 'igSetNextWindowSizeConstraints']
fn set_next_window_size_constraints(size_min ImVec2, size_max ImVec2, custom_callback C.ImGuiSizeCallback, custom_callback_data voidptr)

@[c: 'igSetNextWindowContentSize']
fn set_next_window_content_size(size ImVec2)

@[c: 'igSetNextWindowCollapsed']
fn set_next_window_collapsed(collapsed bool, cond Cond)

@[c: 'igSetNextWindowFocus']
fn set_next_window_focus()

@[c: 'igSetNextWindowScroll']
fn set_next_window_scroll(scroll ImVec2)

@[c: 'igSetNextWindowBgAlpha']
fn set_next_window_bg_alpha(alpha f32)

@[c: 'igSetNextWindowViewport']
fn set_next_window_viewport(viewport_id ID)

@[c: 'igSetWindowPos_Vec2']
fn set_window_pos_vec2(pos ImVec2, cond Cond)

@[c: 'igSetWindowSize_Vec2']
fn set_window_size_vec2(size ImVec2, cond Cond)

@[c: 'igSetWindowCollapsed_Bool']
fn set_window_collapsed_bool(collapsed bool, cond Cond)

@[c: 'igSetWindowFocus_Nil']
fn set_window_focus_nil()

@[c: 'igSetWindowFontScale']
fn set_window_font_scale(scale f32)

@[c: 'igSetWindowPos_Str']
fn set_window_pos_str(name &i8, pos ImVec2, cond Cond)

@[c: 'igSetWindowSize_Str']
fn set_window_size_str(name &i8, size ImVec2, cond Cond)

@[c: 'igSetWindowCollapsed_Str']
fn set_window_collapsed_str(name &i8, collapsed bool, cond Cond)

@[c: 'igSetWindowFocus_Str']
fn set_window_focus_str(name &i8)

@[c: 'igGetScrollX']
fn get_scroll_x() f32

@[c: 'igGetScrollY']
fn get_scroll_y() f32

@[c: 'igSetScrollX_Float']
fn set_scroll_x_float(scroll_x f32)

@[c: 'igSetScrollY_Float']
fn set_scroll_y_float(scroll_y f32)

@[c: 'igGetScrollMaxX']
fn get_scroll_max_x() f32

@[c: 'igGetScrollMaxY']
fn get_scroll_max_y() f32

@[c: 'igSetScrollHereX']
fn set_scroll_here_x(center_x_ratio f32)

@[c: 'igSetScrollHereY']
fn set_scroll_here_y(center_y_ratio f32)

@[c: 'igSetScrollFromPosX_Float']
fn set_scroll_from_pos_x_float(local_x f32, center_x_ratio f32)

@[c: 'igSetScrollFromPosY_Float']
fn set_scroll_from_pos_y_float(local_y f32, center_y_ratio f32)

@[c: 'igPushFont']
fn push_font(font &ImFont)

@[c: 'igPopFont']
fn pop_font()

@[c: 'igPushStyleColor_U32']
fn push_style_color_u32(idx Col, col ImU32)

@[c: 'igPushStyleColor_Vec4']
fn push_style_color_vec4(idx Col, col C.ImVec4)

@[c: 'igPopStyleColor']
fn pop_style_color(count int)

@[c: 'igPushStyleVar_Float']
fn push_style_var_float(idx StyleVar, val f32)

@[c: 'igPushStyleVar_Vec2']
fn push_style_var_vec2(idx StyleVar, val ImVec2)

@[c: 'igPushStyleVarX']
fn push_style_var_x(idx StyleVar, val_x f32)

@[c: 'igPushStyleVarY']
fn push_style_var_y(idx StyleVar, val_y f32)

@[c: 'igPopStyleVar']
fn pop_style_var(count int)

@[c: 'igPushItemFlag']
fn push_item_flag(option ItemFlags, enabled bool)

@[c: 'igPopItemFlag']
fn pop_item_flag()

@[c: 'igPushItemWidth']
fn push_item_width(item_width f32)

@[c: 'igPopItemWidth']
fn pop_item_width()

@[c: 'igSetNextItemWidth']
fn set_next_item_width(item_width f32)

@[c: 'igCalcItemWidth']
fn calc_item_width() f32

@[c: 'igPushTextWrapPos']
fn push_text_wrap_pos(wrap_local_pos_x f32)

@[c: 'igPopTextWrapPos']
fn pop_text_wrap_pos()

@[c: 'igGetFont']
fn get_font() &ImFont

@[c: 'igGetFontSize']
fn get_font_size() f32

@[c: 'igGetFontTexUvWhitePixel']
fn get_font_tex_uv_white_pixel(p_out &ImVec2)

@[c: 'igGetColorU32_Col']
fn get_color_u32_col(idx Col, alpha_mul f32) ImU32

@[c: 'igGetColorU32_Vec4']
fn get_color_u32_vec4(col C.ImVec4) ImU32

@[c: 'igGetColorU32_U32']
fn get_color_u32_u32(col ImU32, alpha_mul f32) ImU32

@[c: 'igGetStyleColorVec4']
fn get_style_color_vec4(idx Col) &C.ImVec4

@[c: 'igGetCursorScreenPos']
fn get_cursor_screen_pos(p_out &ImVec2)

@[c: 'igSetCursorScreenPos']
fn set_cursor_screen_pos(pos ImVec2)

@[c: 'igGetContentRegionAvail']
fn get_content_region_avail(p_out &ImVec2)

@[c: 'igGetCursorPos']
fn get_cursor_pos(p_out &ImVec2)

@[c: 'igGetCursorPosX']
fn get_cursor_pos_x() f32

@[c: 'igGetCursorPosY']
fn get_cursor_pos_y() f32

@[c: 'igSetCursorPos']
fn set_cursor_pos(local_pos ImVec2)

@[c: 'igSetCursorPosX']
fn set_cursor_pos_x(local_x f32)

@[c: 'igSetCursorPosY']
fn set_cursor_pos_y(local_y f32)

@[c: 'igGetCursorStartPos']
fn get_cursor_start_pos(p_out &ImVec2)

@[c: 'igSeparator']
fn separator()

@[c: 'igSameLine']
fn same_line(offset_from_start_x f32, spacing f32)

@[c: 'igNewLine']
fn new_line()

@[c: 'igSpacing']
fn spacing()

@[c: 'igDummy']
fn dummy(size ImVec2)

@[c: 'igIndent']
fn indent(indent_w f32)

@[c: 'igUnindent']
fn unindent(indent_w f32)

@[c: 'igBeginGroup']
fn begin_group()

@[c: 'igEndGroup']
fn end_group()

@[c: 'igAlignTextToFramePadding']
fn align_text_to_frame_padding()

@[c: 'igGetTextLineHeight']
fn get_text_line_height() f32

@[c: 'igGetTextLineHeightWithSpacing']
fn get_text_line_height_with_spacing() f32

@[c: 'igGetFrameHeight']
fn get_frame_height() f32

@[c: 'igGetFrameHeightWithSpacing']
fn get_frame_height_with_spacing() f32

@[c: 'igPushID_Str']
fn push_id_str(str_id &i8)

@[c: 'igPushID_StrStr']
fn push_id_str_str(str_id_begin &i8, str_id_end &i8)

@[c: 'igPushID_Ptr']
fn push_id_ptr(ptr_id voidptr)

@[c: 'igPushID_Int']
fn push_id_int(int_id int)

@[c: 'igPopID']
fn pop_id()

@[c: 'igGetID_Str']
fn get_id_str(str_id &i8) ID

@[c: 'igGetID_StrStr']
fn get_id_str_str(str_id_begin &i8, str_id_end &i8) ID

@[c: 'igGetID_Ptr']
fn get_id_ptr(ptr_id voidptr) ID

@[c: 'igGetID_Int']
fn get_id_int(int_id int) ID

@[c: 'igTextUnformatted']
fn text_unformatted(text &i8, text_end &i8)

@[c: 'igText']
@[c2v_variadic]
fn text(fmt ...&i8)

@[c: 'igTextV']
fn text_v(fmt &i8, args C.va_list)

@[c: 'igTextColored']
@[c2v_variadic]
fn text_colored(col C.ImVec4, fmt ...&i8)

@[c: 'igTextColoredV']
fn text_colored_v(col C.ImVec4, fmt &i8, args C.va_list)

@[c: 'igTextDisabled']
@[c2v_variadic]
fn text_disabled(fmt ...&i8)

@[c: 'igTextDisabledV']
fn text_disabled_v(fmt &i8, args C.va_list)

@[c: 'igTextWrapped']
@[c2v_variadic]
fn text_wrapped(fmt ...&i8)

@[c: 'igTextWrappedV']
fn text_wrapped_v(fmt &i8, args C.va_list)

@[c: 'igLabelText']
@[c2v_variadic]
fn label_text(label &i8, fmt ...&i8)

@[c: 'igLabelTextV']
fn label_text_v(label &i8, fmt &i8, args C.va_list)

@[c: 'igBulletText']
@[c2v_variadic]
fn bullet_text(fmt ...&i8)

@[c: 'igBulletTextV']
fn bullet_text_v(fmt &i8, args C.va_list)

@[c: 'igSeparatorText']
fn separator_text(label &i8)

@[c: 'igButton']
fn button(label &i8, size ImVec2) bool

@[c: 'igSmallButton']
fn small_button(label &i8) bool

@[c: 'igInvisibleButton']
fn invisible_button(str_id &i8, size ImVec2, flags ButtonFlags) bool

@[c: 'igArrowButton']
fn arrow_button(str_id &i8, dir Dir) bool

@[c: 'igCheckbox']
fn checkbox(label &i8, v &bool) bool

@[c: 'igCheckboxFlags_IntPtr']
fn checkbox_flags_int_ptr(label &i8, flags &int, flags_value int) bool

@[c: 'igCheckboxFlags_UintPtr']
fn checkbox_flags_uint_ptr(label &i8, flags &u32, flags_value u32) bool

@[c: 'igRadioButton_Bool']
fn radio_button_bool(label &i8, active bool) bool

@[c: 'igRadioButton_IntPtr']
fn radio_button_int_ptr(label &i8, v &int, v_button int) bool

@[c: 'igProgressBar']
fn progress_bar(fraction f32, size_arg ImVec2, overlay &i8)

@[c: 'igBullet']
fn bullet()

@[c: 'igTextLink']
fn text_link(label &i8) bool

@[c: 'igTextLinkOpenURL']
fn text_link_open_url(label &i8, url &i8)

@[c: 'igImage']
fn image(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2)

@[c: 'igImageWithBg']
fn image_with_bg(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col C.ImVec4, tint_col C.ImVec4)

@[c: 'igImageButton']
fn image_button(str_id &i8, user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col C.ImVec4, tint_col C.ImVec4) bool

@[c: 'igBeginCombo']
fn begin_combo(label &i8, preview_value &i8, flags ComboFlags) bool

@[c: 'igEndCombo']
fn end_combo()

@[c: 'igCombo_Str_arr']
fn combo_str_arr(label &i8, current_item &int, items &&u8, items_count int, popup_max_height_in_items int) bool

@[c: 'igCombo_Str']
fn combo_str(label &i8, current_item &int, items_separated_by_zeros &i8, popup_max_height_in_items int) bool

@[c: 'igCombo_FnStrPtr']
fn combo_fn_str_ptr(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int, popup_max_height_in_items int) bool

@[c: 'igDragFloat']
fn drag_float(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloat2']
fn drag_float2(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloat3']
fn drag_float3(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloat4']
fn drag_float4(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloatRange2']
fn drag_float_range2(label &i8, v_current_min &f32, v_current_max &f32, v_speed f32, v_min f32, v_max f32, format &i8, format_max &i8, flags SliderFlags) bool

@[c: 'igDragInt']
fn drag_int(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragInt2']
fn drag_int2(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragInt3']
fn drag_int3(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragInt4']
fn drag_int4(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragIntRange2']
fn drag_int_range2(label &i8, v_current_min &int, v_current_max &int, v_speed f32, v_min int, v_max int, format &i8, format_max &i8, flags SliderFlags) bool

@[c: 'igDragScalar']
fn drag_scalar(label &i8, data_type DataType, p_data voidptr, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igDragScalarN']
fn drag_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat']
fn slider_float(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat2']
fn slider_float2(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat3']
fn slider_float3(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat4']
fn slider_float4(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderAngle']
fn slider_angle(label &i8, v_rad &f32, v_degrees_min f32, v_degrees_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt']
fn slider_int(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt2']
fn slider_int2(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt3']
fn slider_int3(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt4']
fn slider_int4(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderScalar']
fn slider_scalar(label &i8, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igSliderScalarN']
fn slider_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igVSliderFloat']
fn vs_lider_float(label &i8, size ImVec2, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igVSliderInt']
fn vs_lider_int(label &i8, size ImVec2, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igVSliderScalar']
fn vs_lider_scalar(label &i8, size ImVec2, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igInputText']
fn input_text(label &i8, buf &i8, buf_size usize, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c: 'igInputTextMultiline']
fn input_text_multiline(label &i8, buf &i8, buf_size usize, size ImVec2, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c: 'igInputTextWithHint']
fn input_text_with_hint(label &i8, hint &i8, buf &i8, buf_size usize, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c: 'igInputFloat']
fn input_float(label &i8, v &f32, step f32, step_fast f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputFloat2']
fn input_float2(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputFloat3']
fn input_float3(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputFloat4']
fn input_float4(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputInt']
fn input_int(label &i8, v &int, step int, step_fast int, flags InputTextFlags) bool

@[c: 'igInputInt2']
fn input_int2(label &i8, v &int, flags InputTextFlags) bool

@[c: 'igInputInt3']
fn input_int3(label &i8, v &int, flags InputTextFlags) bool

@[c: 'igInputInt4']
fn input_int4(label &i8, v &int, flags InputTextFlags) bool

@[c: 'igInputDouble']
fn input_double(label &i8, v &f64, step f64, step_fast f64, format &i8, flags InputTextFlags) bool

@[c: 'igInputScalar']
fn input_scalar(label &i8, data_type DataType, p_data voidptr, p_step voidptr, p_step_fast voidptr, format &i8, flags InputTextFlags) bool

@[c: 'igInputScalarN']
fn input_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, p_step voidptr, p_step_fast voidptr, format &i8, flags InputTextFlags) bool

@[c: 'igColorEdit3']
fn color_edit3(label &i8, col &f32, flags ColorEditFlags) bool

@[c: 'igColorEdit4']
fn color_edit4(label &i8, col &f32, flags ColorEditFlags) bool

@[c: 'igColorPicker3']
fn color_picker3(label &i8, col &f32, flags ColorEditFlags) bool

@[c: 'igColorPicker4']
fn color_picker4(label &i8, col &f32, flags ColorEditFlags, ref_col &f32) bool

@[c: 'igColorButton']
fn color_button(desc_id &i8, col C.ImVec4, flags ColorEditFlags, size ImVec2) bool

@[c: 'igSetColorEditOptions']
fn set_color_edit_options(flags ColorEditFlags)

@[c: 'igTreeNode_Str']
fn tree_node_str(label &i8) bool

@[c: 'igTreeNode_StrStr']
@[c2v_variadic]
fn tree_node_str_str(str_id &i8, fmt ...&i8) bool

@[c: 'igTreeNode_Ptr']
@[c2v_variadic]
fn tree_node_ptr(ptr_id voidptr, fmt ...&i8) bool

@[c: 'igTreeNodeV_Str']
fn tree_node_v_str(str_id &i8, fmt &i8, args C.va_list) bool

@[c: 'igTreeNodeV_Ptr']
fn tree_node_v_ptr(ptr_id voidptr, fmt &i8, args C.va_list) bool

@[c: 'igTreeNodeEx_Str']
fn tree_node_ex_str(label &i8, flags TreeNodeFlags) bool

@[c: 'igTreeNodeEx_StrStr']
@[c2v_variadic]
fn tree_node_ex_str_str(str_id &i8, flags TreeNodeFlags, fmt ...&i8) bool

@[c: 'igTreeNodeEx_Ptr']
@[c2v_variadic]
fn tree_node_ex_ptr(ptr_id voidptr, flags TreeNodeFlags, fmt ...&i8) bool

@[c: 'igTreeNodeExV_Str']
fn tree_node_ex_v_str(str_id &i8, flags TreeNodeFlags, fmt &i8, args C.va_list) bool

@[c: 'igTreeNodeExV_Ptr']
fn tree_node_ex_v_ptr(ptr_id voidptr, flags TreeNodeFlags, fmt &i8, args C.va_list) bool

@[c: 'igTreePush_Str']
fn tree_push_str(str_id &i8)

@[c: 'igTreePush_Ptr']
fn tree_push_ptr(ptr_id voidptr)

@[c: 'igTreePop']
fn tree_pop()

@[c: 'igGetTreeNodeToLabelSpacing']
fn get_tree_node_to_label_spacing() f32

@[c: 'igCollapsingHeader_TreeNodeFlags']
fn collapsing_header_tree_node_flags(label &i8, flags TreeNodeFlags) bool

@[c: 'igCollapsingHeader_BoolPtr']
fn collapsing_header_bool_ptr(label &i8, p_visible &bool, flags TreeNodeFlags) bool

@[c: 'igSetNextItemOpen']
fn set_next_item_open(is_open bool, cond Cond)

@[c: 'igSetNextItemStorageID']
fn set_next_item_storage_id(storage_id ID)

@[c: 'igSelectable_Bool']
fn selectable_bool(label &i8, selected bool, flags SelectableFlags, size ImVec2) bool

@[c: 'igSelectable_BoolPtr']
fn selectable_bool_ptr(label &i8, p_selected &bool, flags SelectableFlags, size ImVec2) bool

@[c: 'igBeginMultiSelect']
fn begin_multi_select(flags MultiSelectFlags, selection_size int, items_count int) &MultiSelectIO

@[c: 'igEndMultiSelect']
fn end_multi_select() &MultiSelectIO

@[c: 'igSetNextItemSelectionUserData']
fn set_next_item_selection_user_data(selection_user_data SelectionUserData)

@[c: 'igIsItemToggledSelection']
fn is_item_toggled_selection() bool

@[c: 'igBeginListBox']
fn begin_list_box(label &i8, size ImVec2) bool

@[c: 'igEndListBox']
fn end_list_box()

@[c: 'igListBox_Str_arr']
fn list_box_str_arr(label &i8, current_item &int, items &&u8, items_count int, height_in_items int) bool

@[c: 'igListBox_FnStrPtr']
fn list_box_fn_str_ptr(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int, height_in_items int) bool

@[c: 'igPlotLines_FloatPtr']
fn plot_lines_float_ptr(label &i8, values &f32, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2, stride int)

@[c: 'igPlotLines_FnFloatPtr']
fn plot_lines_fn_float_ptr(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2)

@[c: 'igPlotHistogram_FloatPtr']
fn plot_histogram_float_ptr(label &i8, values &f32, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2, stride int)

@[c: 'igPlotHistogram_FnFloatPtr']
fn plot_histogram_fn_float_ptr(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2)

@[c: 'igValue_Bool']
fn value_bool(prefix &i8, b bool)

@[c: 'igValue_Int']
fn value_int(prefix &i8, v int)

@[c: 'igValue_Uint']
fn value_uint(prefix &i8, v u32)

@[c: 'igValue_Float']
fn value_float(prefix &i8, v f32, float_format &i8)

@[c: 'igBeginMenuBar']
fn begin_menu_bar() bool

@[c: 'igEndMenuBar']
fn end_menu_bar()

@[c: 'igBeginMainMenuBar']
fn begin_main_menu_bar() bool

@[c: 'igEndMainMenuBar']
fn end_main_menu_bar()

@[c: 'igBeginMenu']
fn begin_menu(label &i8, enabled bool) bool

@[c: 'igEndMenu']
fn end_menu()

@[c: 'igMenuItem_Bool']
fn menu_item_bool(label &i8, shortcut &i8, selected bool, enabled bool) bool

@[c: 'igMenuItem_BoolPtr']
fn menu_item_bool_ptr(label &i8, shortcut &i8, p_selected &bool, enabled bool) bool

@[c: 'igBeginTooltip']
fn begin_tooltip() bool

@[c: 'igEndTooltip']
fn end_tooltip()

@[c: 'igSetTooltip']
@[c2v_variadic]
fn set_tooltip(fmt ...&i8)

@[c: 'igSetTooltipV']
fn set_tooltip_v(fmt &i8, args C.va_list)

@[c: 'igBeginItemTooltip']
fn begin_item_tooltip() bool

@[c: 'igSetItemTooltip']
@[c2v_variadic]
fn set_item_tooltip(fmt ...&i8)

@[c: 'igSetItemTooltipV']
fn set_item_tooltip_v(fmt &i8, args C.va_list)

@[c: 'igBeginPopup']
fn begin_popup(str_id &i8, flags WindowFlags) bool

@[c: 'igBeginPopupModal']
fn begin_popup_modal(name &i8, p_open &bool, flags WindowFlags) bool

@[c: 'igEndPopup']
fn end_popup()

@[c: 'igOpenPopup_Str']
fn open_popup_str(str_id &i8, popup_flags PopupFlags)

@[c: 'igOpenPopup_ID']
fn open_popup_id(id ID, popup_flags PopupFlags)

@[c: 'igOpenPopupOnItemClick']
fn open_popup_on_item_click(str_id &i8, popup_flags PopupFlags)

@[c: 'igCloseCurrentPopup']
fn close_current_popup()

@[c: 'igBeginPopupContextItem']
fn begin_popup_context_item(str_id &i8, popup_flags PopupFlags) bool

@[c: 'igBeginPopupContextWindow']
fn begin_popup_context_window(str_id &i8, popup_flags PopupFlags) bool

@[c: 'igBeginPopupContextVoid']
fn begin_popup_context_void(str_id &i8, popup_flags PopupFlags) bool

@[c: 'igIsPopupOpen_Str']
fn is_popup_open_str(str_id &i8, flags PopupFlags) bool

@[c: 'igBeginTable']
fn begin_table(str_id &i8, columns int, flags TableFlags, outer_size ImVec2, inner_width f32) bool

@[c: 'igEndTable']
fn end_table()

@[c: 'igTableNextRow']
fn table_next_row(row_flags TableRowFlags, min_row_height f32)

@[c: 'igTableNextColumn']
fn table_next_column() bool

@[c: 'igTableSetColumnIndex']
fn table_set_column_index(column_n int) bool

@[c: 'igTableSetupColumn']
fn table_setup_column(label &i8, flags TableColumnFlags, init_width_or_weight f32, user_id ID)

@[c: 'igTableSetupScrollFreeze']
fn table_setup_scroll_freeze(cols int, rows int)

@[c: 'igTableHeader']
fn table_header(label &i8)

@[c: 'igTableHeadersRow']
fn table_headers_row()

@[c: 'igTableAngledHeadersRow']
fn table_angled_headers_row()

@[c: 'igTableGetSortSpecs']
fn table_get_sort_specs() &TableSortSpecs

@[c: 'igTableGetColumnCount']
fn table_get_column_count() int

@[c: 'igTableGetColumnIndex']
fn table_get_column_index() int

@[c: 'igTableGetRowIndex']
fn table_get_row_index() int

@[c: 'igTableGetColumnName_Int']
fn table_get_column_name_int(column_n int) &i8

@[c: 'igTableGetColumnFlags']
fn table_get_column_flags(column_n int) TableColumnFlags

@[c: 'igTableSetColumnEnabled']
fn table_set_column_enabled(column_n int, v bool)

@[c: 'igTableGetHoveredColumn']
fn table_get_hovered_column() int

@[c: 'igTableSetBgColor']
fn table_set_bg_color(target TableBgTarget, color ImU32, column_n int)

@[c: 'igColumns']
fn columns(count int, id &i8, borders bool)

@[c: 'igNextColumn']
fn next_column()

@[c: 'igGetColumnIndex']
fn get_column_index() int

@[c: 'igGetColumnWidth']
fn get_column_width(column_index int) f32

@[c: 'igSetColumnWidth']
fn set_column_width(column_index int, width f32)

@[c: 'igGetColumnOffset']
fn get_column_offset(column_index int) f32

@[c: 'igSetColumnOffset']
fn set_column_offset(column_index int, offset_x f32)

@[c: 'igGetColumnsCount']
fn get_columns_count() int

@[c: 'igBeginTabBar']
fn begin_tab_bar(str_id &i8, flags ImGuiTabBarFlags) bool

@[c: 'igEndTabBar']
fn end_tab_bar()

@[c: 'igBeginTabItem']
fn begin_tab_item(label &i8, p_open &bool, flags TabItemFlags) bool

@[c: 'igEndTabItem']
fn end_tab_item()

@[c: 'igTabItemButton']
fn tab_item_button(label &i8, flags TabItemFlags) bool

@[c: 'igSetTabItemClosed']
fn set_tab_item_closed(tab_or_docked_window_label &i8)

@[c: 'igDockSpace']
fn dock_space(dockspace_id ID, size ImVec2, flags DockNodeFlags, window_class &WindowClass) ID

@[c: 'igDockSpaceOverViewport']
fn dock_space_over_viewport(dockspace_id ID, viewport &Viewport, flags DockNodeFlags, window_class &WindowClass) ID

@[c: 'igSetNextWindowDockID']
fn set_next_window_dock_id(dock_id ID, cond Cond)

@[c: 'igSetNextWindowClass']
fn set_next_window_class(window_class &WindowClass)

@[c: 'igGetWindowDockID']
fn get_window_dock_id() ID

@[c: 'igIsWindowDocked']
fn is_window_docked() bool

@[c: 'igLogToTTY']
fn log_to_tty(auto_open_depth int)

@[c: 'igLogToFile']
fn log_to_file(auto_open_depth int, filename &i8)

@[c: 'igLogToClipboard']
fn log_to_clipboard(auto_open_depth int)

@[c: 'igLogFinish']
fn log_finish()

@[c: 'igLogButtons']
fn log_buttons()

@[c: 'igLogTextV']
fn log_text_v(fmt &i8, args C.va_list)

@[c: 'igBeginDragDropSource']
fn begin_drag_drop_source(flags DragDropFlags) bool

@[c: 'igSetDragDropPayload']
fn set_drag_drop_payload(type_ &i8, data voidptr, sz usize, cond Cond) bool

@[c: 'igEndDragDropSource']
fn end_drag_drop_source()

@[c: 'igBeginDragDropTarget']
fn begin_drag_drop_target() bool

@[c: 'igAcceptDragDropPayload']
fn accept_drag_drop_payload(type_ &i8, flags DragDropFlags) &Payload

@[c: 'igEndDragDropTarget']
fn end_drag_drop_target()

@[c: 'igGetDragDropPayload']
fn get_drag_drop_payload() &Payload

@[c: 'igBeginDisabled']
fn begin_disabled(disabled bool)

@[c: 'igEndDisabled']
fn end_disabled()

@[c: 'igPushClipRect']
fn push_clip_rect(clip_rect_min ImVec2, clip_rect_max ImVec2, intersect_with_current_clip_rect bool)

@[c: 'igPopClipRect']
fn pop_clip_rect()

@[c: 'igSetItemDefaultFocus']
fn set_item_default_focus()

@[c: 'igSetKeyboardFocusHere']
fn set_keyboard_focus_here(offset int)

@[c: 'igSetNavCursorVisible']
fn set_nav_cursor_visible(visible bool)

@[c: 'igSetNextItemAllowOverlap']
fn set_next_item_allow_overlap()

@[c: 'igIsItemHovered']
fn is_item_hovered(flags HoveredFlags) bool

@[c: 'igIsItemActive']
fn is_item_active() bool

@[c: 'igIsItemFocused']
fn is_item_focused() bool

@[c: 'igIsItemClicked']
fn is_item_clicked(mouse_button MouseButton) bool

@[c: 'igIsItemVisible']
fn is_item_visible() bool

@[c: 'igIsItemEdited']
fn is_item_edited() bool

@[c: 'igIsItemActivated']
fn is_item_activated() bool

@[c: 'igIsItemDeactivated']
fn is_item_deactivated() bool

@[c: 'igIsItemDeactivatedAfterEdit']
fn is_item_deactivated_after_edit() bool

@[c: 'igIsItemToggledOpen']
fn is_item_toggled_open() bool

@[c: 'igIsAnyItemHovered']
fn is_any_item_hovered() bool

@[c: 'igIsAnyItemActive']
fn is_any_item_active() bool

@[c: 'igIsAnyItemFocused']
fn is_any_item_focused() bool

@[c: 'igGetItemID']
fn get_item_id() ID

@[c: 'igGetItemRectMin']
fn get_item_rect_min(p_out &ImVec2)

@[c: 'igGetItemRectMax']
fn get_item_rect_max(p_out &ImVec2)

@[c: 'igGetItemRectSize']
fn get_item_rect_size(p_out &ImVec2)

@[c: 'igGetMainViewport']
fn get_main_viewport() &Viewport

@[c: 'igGetBackgroundDrawList']
fn get_background_draw_list(viewport &Viewport) &ImDrawList

@[c: 'igGetForegroundDrawList_ViewportPtr']
fn get_foreground_draw_list_viewport_ptr(viewport &Viewport) &ImDrawList

@[c: 'igIsRectVisible_Nil']
fn is_rect_visible_nil(size ImVec2) bool

@[c: 'igIsRectVisible_Vec2']
fn is_rect_visible_vec2(rect_min ImVec2, rect_max ImVec2) bool

@[c: 'igGetTime']
fn get_time() f64

@[c: 'igGetFrameCount']
fn get_frame_count() int

@[c: 'igGetDrawListSharedData']
fn get_draw_list_shared_data() &ImDrawListSharedData

@[c: 'igGetStyleColorName']
fn get_style_color_name(idx Col) &i8

@[c: 'igSetStateStorage']
fn set_state_storage(storage &Storage)

@[c: 'igGetStateStorage']
fn get_state_storage() &Storage

@[c: 'igCalcTextSize']
fn calc_text_size(p_out &ImVec2, text &i8, text_end &i8, hide_text_after_double_hash bool, wrap_width f32)

@[c: 'igColorConvertU32ToFloat4']
fn color_convert_u32_to_float4(p_out &C.ImVec4, in_ ImU32)

@[c: 'igColorConvertFloat4ToU32']
fn color_convert_float4_to_u32(in_ C.ImVec4) ImU32

@[c: 'igColorConvertRGBtoHSV']
fn color_convert_rgb_to_hsv(r f32, g f32, b f32, out_h &f32, out_s &f32, out_v &f32)

@[c: 'igColorConvertHSVtoRGB']
fn color_convert_hsv_to_rgb(h f32, s f32, v f32, out_r &f32, out_g &f32, out_b &f32)

@[c: 'igIsKeyDown_Nil']
fn is_key_down_nil(key Key) bool

@[c: 'igIsKeyPressed_Bool']
fn is_key_pressed_bool(key Key, repeat bool) bool

@[c: 'igIsKeyReleased_Nil']
fn is_key_released_nil(key Key) bool

@[c: 'igIsKeyChordPressed_Nil']
fn is_key_chord_pressed_nil(key_chord KeyChord) bool

@[c: 'igGetKeyPressedAmount']
fn get_key_pressed_amount(key Key, repeat_delay f32, rate f32) int

@[c: 'igGetKeyName']
fn get_key_name(key Key) &i8

@[c: 'igSetNextFrameWantCaptureKeyboard']
fn set_next_frame_want_capture_keyboard(want_capture_keyboard bool)

@[c: 'igShortcut_Nil']
fn shortcut_nil(key_chord KeyChord, flags InputFlags) bool

@[c: 'igSetNextItemShortcut']
fn set_next_item_shortcut(key_chord KeyChord, flags InputFlags)

@[c: 'igSetItemKeyOwner_Nil']
fn set_item_key_owner_nil(key Key)

@[c: 'igIsMouseDown_Nil']
fn is_mouse_down_nil(button MouseButton) bool

@[c: 'igIsMouseClicked_Bool']
fn is_mouse_clicked_bool(button MouseButton, repeat bool) bool

@[c: 'igIsMouseReleased_Nil']
fn is_mouse_released_nil(button MouseButton) bool

@[c: 'igIsMouseDoubleClicked_Nil']
fn is_mouse_double_clicked_nil(button MouseButton) bool

@[c: 'igIsMouseReleasedWithDelay']
fn is_mouse_released_with_delay(button MouseButton, delay f32) bool

@[c: 'igGetMouseClickedCount']
fn get_mouse_clicked_count(button MouseButton) int

@[c: 'igIsMouseHoveringRect']
fn is_mouse_hovering_rect(r_min ImVec2, r_max ImVec2, clip bool) bool

@[c: 'igIsMousePosValid']
fn is_mouse_pos_valid(mouse_pos &ImVec2) bool

@[c: 'igIsAnyMouseDown']
fn is_any_mouse_down() bool

@[c: 'igGetMousePos']
fn get_mouse_pos(p_out &ImVec2)

@[c: 'igGetMousePosOnOpeningCurrentPopup']
fn get_mouse_pos_on_opening_current_popup(p_out &ImVec2)

@[c: 'igIsMouseDragging']
fn is_mouse_dragging(button MouseButton, lock_threshold f32) bool

@[c: 'igGetMouseDragDelta']
fn get_mouse_drag_delta(p_out &ImVec2, button MouseButton, lock_threshold f32)

@[c: 'igResetMouseDragDelta']
fn reset_mouse_drag_delta(button MouseButton)

@[c: 'igGetMouseCursor']
fn get_mouse_cursor() MouseCursor

@[c: 'igSetMouseCursor']
fn set_mouse_cursor(cursor_type MouseCursor)

@[c: 'igSetNextFrameWantCaptureMouse']
fn set_next_frame_want_capture_mouse(want_capture_mouse bool)

@[c: 'igGetClipboardText']
fn get_clipboard_text() &i8

@[c: 'igSetClipboardText']
fn set_clipboard_text(text &i8)

@[c: 'igLoadIniSettingsFromDisk']
fn load_ini_settings_from_disk(ini_filename &i8)

@[c: 'igLoadIniSettingsFromMemory']
fn load_ini_settings_from_memory(ini_data &i8, ini_size usize)

@[c: 'igSaveIniSettingsToDisk']
fn save_ini_settings_to_disk(ini_filename &i8)

@[c: 'igSaveIniSettingsToMemory']
fn save_ini_settings_to_memory(out_ini_size &usize) &i8

@[c: 'igDebugTextEncoding']
fn debug_text_encoding(text &i8)

@[c: 'igDebugFlashStyleColor']
fn debug_flash_style_color(idx Col)

@[c: 'igDebugStartItemPicker']
fn debug_start_item_picker()

@[c: 'igDebugCheckVersionAndDataLayout']
fn debug_check_version_and_data_layout(version_str &i8, sz_io usize, sz_style usize, sz_vec2 usize, sz_vec4 usize, sz_drawvert usize, sz_drawidx usize) bool

@[c: 'igDebugLog']
@[c2v_variadic]
fn debug_log(fmt ...&i8)

@[c: 'igDebugLogV']
fn debug_log_v(fmt &i8, args C.va_list)

@[c: 'igSetAllocatorFunctions']
fn set_allocator_functions(alloc_func MemAllocFunc, free_func MemFreeFunc, user_data voidptr)

@[c: 'igGetAllocatorFunctions']
fn get_allocator_functions(p_alloc_func &MemAllocFunc, p_free_func &MemFreeFunc, p_user_data &voidptr)

@[c: 'igMemAlloc']
fn mem_alloc(size usize) voidptr

@[c: 'igMemFree']
fn mem_free(ptr voidptr)

@[c: 'igUpdatePlatformWindows']
fn update_platform_windows()

@[c: 'igRenderPlatformWindowsDefault']
fn render_platform_windows_default(platform_render_arg voidptr, renderer_render_arg voidptr)

@[c: 'igDestroyPlatformWindows']
fn destroy_platform_windows()

@[c: 'igFindViewportByID']
fn find_viewport_by_id(id ID) &Viewport

@[c: 'igFindViewportByPlatformHandle']
fn find_viewport_by_platform_handle(platform_handle voidptr) &Viewport

@[c: 'ImGuiTableSortSpecs_ImGuiTableSortSpecs']
fn table_sort_specs_im_gui_table_sort_specs() &TableSortSpecs

@[c: 'ImGuiTableSortSpecs_ImGuiTableSortSpecs_Construct']
fn table_sort_specs_im_gui_table_sort_specs_construct(self &TableSortSpecs)

@[c: 'ImGuiTableSortSpecs_destroy']
fn table_sort_specs_destroy(self &TableSortSpecs)

@[c: 'ImGuiTableColumnSortSpecs_ImGuiTableColumnSortSpecs']
fn table_column_sort_specs_im_gui_table_column_sort_specs() &TableColumnSortSpecs

@[c: 'ImGuiTableColumnSortSpecs_ImGuiTableColumnSortSpecs_Construct']
fn table_column_sort_specs_im_gui_table_column_sort_specs_construct(self &TableColumnSortSpecs)

@[c: 'ImGuiTableColumnSortSpecs_destroy']
fn table_column_sort_specs_destroy(self &TableColumnSortSpecs)

@[c: 'ImGuiStyle_ImGuiStyle']
fn style_im_gui_style() &Style

@[c: 'ImGuiStyle_ImGuiStyle_Construct']
fn style_im_gui_style_construct(self &Style)

@[c: 'ImGuiStyle_destroy']
fn style_destroy(self &Style)

@[c: 'ImGuiStyle_ScaleAllSizes']
fn style_scale_all_sizes(self &Style, scale_factor f32)

@[c: 'ImGuiIO_AddKeyEvent']
fn io_add_key_event(self &IO, key Key, down bool)

@[c: 'ImGuiIO_AddKeyAnalogEvent']
fn io_add_key_analog_event(self &IO, key Key, down bool, v f32)

@[c: 'ImGuiIO_AddMousePosEvent']
fn io_add_mouse_pos_event(self &IO, x f32, y f32)

@[c: 'ImGuiIO_AddMouseButtonEvent']
fn io_add_mouse_button_event(self &IO, button int, down bool)

@[c: 'ImGuiIO_AddMouseWheelEvent']
fn io_add_mouse_wheel_event(self &IO, wheel_x f32, wheel_y f32)

@[c: 'ImGuiIO_AddMouseSourceEvent']
fn io_add_mouse_source_event(self &IO, source MouseSource)

@[c: 'ImGuiIO_AddMouseViewportEvent']
fn io_add_mouse_viewport_event(self &IO, id ID)

@[c: 'ImGuiIO_AddFocusEvent']
fn io_add_focus_event(self &IO, focused bool)

@[c: 'ImGuiIO_AddInputCharacter']
fn io_add_input_character(self &IO, c u32)

@[c: 'ImGuiIO_AddInputCharacterUTF16']
fn io_add_input_character_utf_16(self &IO, c ImWchar16)

@[c: 'ImGuiIO_AddInputCharactersUTF8']
fn io_add_input_characters_utf_8(self &IO, str &i8)

@[c: 'ImGuiIO_SetKeyEventNativeData']
fn io_set_key_event_native_data(self &IO, key Key, native_keycode int, native_scancode int, native_legacy_index int)

@[c: 'ImGuiIO_SetAppAcceptingEvents']
fn io_set_app_accepting_events(self &IO, accepting_events bool)

@[c: 'ImGuiIO_ClearEventsQueue']
fn io_clear_events_queue(self &IO)

@[c: 'ImGuiIO_ClearInputKeys']
fn io_clear_input_keys(self &IO)

@[c: 'ImGuiIO_ClearInputMouse']
fn io_clear_input_mouse(self &IO)

@[c: 'ImGuiIO_ImGuiIO']
fn io_im_gui_io() &IO

@[c: 'ImGuiIO_ImGuiIO_Construct']
fn io_im_gui_io_construct(self &IO)

@[c: 'ImGuiIO_destroy']
fn io_destroy(self &IO)

@[c: 'ImGuiInputTextCallbackData_ImGuiInputTextCallbackData']
fn input_text_callback_data_im_gui_input_text_callback_data() &ImGuiInputTextCallbackData

@[c: 'ImGuiInputTextCallbackData_ImGuiInputTextCallbackData_Construct']
fn input_text_callback_data_im_gui_input_text_callback_data_construct(self &ImGuiInputTextCallbackData)

@[c: 'ImGuiInputTextCallbackData_destroy']
fn input_text_callback_data_destroy(self &ImGuiInputTextCallbackData)

@[c: 'ImGuiInputTextCallbackData_DeleteChars']
fn input_text_callback_data_delete_chars(self &ImGuiInputTextCallbackData, pos int, bytes_count int)

@[c: 'ImGuiInputTextCallbackData_InsertChars']
fn input_text_callback_data_insert_chars(self &ImGuiInputTextCallbackData, pos int, text &i8, text_end &i8)

@[c: 'ImGuiInputTextCallbackData_SelectAll']
fn input_text_callback_data_select_all(self &ImGuiInputTextCallbackData)

@[c: 'ImGuiInputTextCallbackData_ClearSelection']
fn input_text_callback_data_clear_selection(self &ImGuiInputTextCallbackData)

@[c: 'ImGuiInputTextCallbackData_HasSelection']
fn input_text_callback_data_has_selection(self &ImGuiInputTextCallbackData) bool

@[c: 'ImGuiWindowClass_ImGuiWindowClass']
fn window_class_im_gui_window_class() &WindowClass

@[c: 'ImGuiWindowClass_ImGuiWindowClass_Construct']
fn window_class_im_gui_window_class_construct(self &WindowClass)

@[c: 'ImGuiWindowClass_destroy']
fn window_class_destroy(self &WindowClass)

@[c: 'ImGuiPayload_ImGuiPayload']
fn payload_im_gui_payload() &Payload

@[c: 'ImGuiPayload_ImGuiPayload_Construct']
fn payload_im_gui_payload_construct(self &Payload)

@[c: 'ImGuiPayload_destroy']
fn payload_destroy(self &Payload)

@[c: 'ImGuiPayload_Clear']
fn payload_clear(self &Payload)

@[c: 'ImGuiPayload_IsDataType']
fn payload_is_data_type(self &Payload, type_ &i8) bool

@[c: 'ImGuiPayload_IsPreview']
fn payload_is_preview(self &Payload) bool

@[c: 'ImGuiPayload_IsDelivery']
fn payload_is_delivery(self &Payload) bool

@[c: 'ImGuiOnceUponAFrame_ImGuiOnceUponAFrame']
fn once_upon_af_rame_im_gui_once_upon_af_rame() &OnceUponAFrame

@[c: 'ImGuiOnceUponAFrame_ImGuiOnceUponAFrame_Construct']
fn once_upon_af_rame_im_gui_once_upon_af_rame_construct(self &OnceUponAFrame)

@[c: 'ImGuiOnceUponAFrame_destroy']
fn once_upon_af_rame_destroy(self &OnceUponAFrame)

@[c: 'ImGuiTextFilter_ImGuiTextFilter']
fn text_filter_im_gui_text_filter(default_filter &i8) &C.ImGuiTextFilter

@[c: 'ImGuiTextFilter_ImGuiTextFilter_Construct']
fn text_filter_im_gui_text_filter_construct(self &C.ImGuiTextFilter, default_filter &i8)

@[c: 'ImGuiTextFilter_destroy']
fn text_filter_destroy(self &C.ImGuiTextFilter)

@[c: 'ImGuiTextFilter_Draw']
fn text_filter_draw(self &C.ImGuiTextFilter, label &i8, width f32) bool

@[c: 'ImGuiTextFilter_PassFilter']
fn text_filter_pass_filter(self &C.ImGuiTextFilter, text &i8, text_end &i8) bool

@[c: 'ImGuiTextFilter_Build']
fn text_filter_build(self &C.ImGuiTextFilter)

@[c: 'ImGuiTextFilter_Clear']
fn text_filter_clear(self &C.ImGuiTextFilter)

@[c: 'ImGuiTextFilter_IsActive']
fn text_filter_is_active(self &C.ImGuiTextFilter) bool

@[c: 'ImGuiTextRange_ImGuiTextRange_Nil']
fn text_range_im_gui_text_range_nil() &TextRange

@[c: 'ImGuiTextRange_ImGuiTextRange_Nil_Construct']
fn text_range_im_gui_text_range_nil_construct(self &TextRange)

@[c: 'ImGuiTextRange_destroy']
fn text_range_destroy(self &TextRange)

@[c: 'ImGuiTextRange_ImGuiTextRange_Str']
fn text_range_im_gui_text_range_str(_b &i8, _e &i8) &TextRange

@[c: 'ImGuiTextRange_ImGuiTextRange_Str_Construct']
fn text_range_im_gui_text_range_str_construct(self &TextRange, _b &i8, _e &i8)

@[c: 'ImGuiTextRange_empty']
fn text_range_empty(self &TextRange) bool

@[c: 'ImGuiTextRange_split']
fn text_range_split(self &TextRange, separator i8, out &ImVector_ImGuiTextRange)

@[c: 'ImGuiTextBuffer_ImGuiTextBuffer']
fn text_buffer_im_gui_text_buffer() &TextBuffer

@[c: 'ImGuiTextBuffer_ImGuiTextBuffer_Construct']
fn text_buffer_im_gui_text_buffer_construct(self &TextBuffer)

@[c: 'ImGuiTextBuffer_destroy']
fn text_buffer_destroy(self &TextBuffer)

@[c: 'ImGuiTextBuffer_begin']
fn text_buffer_begin(self &TextBuffer) &i8

@[c: 'ImGuiTextBuffer_end']
fn text_buffer_end(self &TextBuffer) &i8

@[c: 'ImGuiTextBuffer_size']
fn text_buffer_size(self &TextBuffer) int

@[c: 'ImGuiTextBuffer_empty']
fn text_buffer_empty(self &TextBuffer) bool

@[c: 'ImGuiTextBuffer_clear']
fn text_buffer_clear(self &TextBuffer)

@[c: 'ImGuiTextBuffer_resize']
fn text_buffer_resize(self &TextBuffer, size int)

@[c: 'ImGuiTextBuffer_reserve']
fn text_buffer_reserve(self &TextBuffer, capacity int)

@[c: 'ImGuiTextBuffer_c_str']
fn text_buffer_c_str(self &TextBuffer) &i8

@[c: 'ImGuiTextBuffer_append']
fn text_buffer_append(self &TextBuffer, str &i8, str_end &i8)

@[c: 'ImGuiTextBuffer_appendfv']
fn text_buffer_appendfv(self &TextBuffer, fmt &i8, args C.va_list)

@[c: 'ImGuiStoragePair_ImGuiStoragePair_Int']
fn storage_pair_im_gui_storage_pair_int(_key ID, _val int) &StoragePair

@[c: 'ImGuiStoragePair_ImGuiStoragePair_Int_Construct']
fn storage_pair_im_gui_storage_pair_int_construct(self &StoragePair, _key ID, _val int)

@[c: 'ImGuiStoragePair_destroy']
fn storage_pair_destroy(self &StoragePair)

@[c: 'ImGuiStoragePair_ImGuiStoragePair_Float']
fn storage_pair_im_gui_storage_pair_float(_key ID, _val f32) &StoragePair

@[c: 'ImGuiStoragePair_ImGuiStoragePair_Float_Construct']
fn storage_pair_im_gui_storage_pair_float_construct(self &StoragePair, _key ID, _val f32)

@[c: 'ImGuiStoragePair_ImGuiStoragePair_Ptr']
fn storage_pair_im_gui_storage_pair_ptr(_key ID, _val voidptr) &StoragePair

@[c: 'ImGuiStoragePair_ImGuiStoragePair_Ptr_Construct']
fn storage_pair_im_gui_storage_pair_ptr_construct(self &StoragePair, _key ID, _val voidptr)

@[c: 'ImGuiStorage_Clear']
fn storage_clear(self &Storage)

@[c: 'ImGuiStorage_GetInt']
fn storage_get_int(self &Storage, key ID, default_val int) int

@[c: 'ImGuiStorage_SetInt']
fn storage_set_int(self &Storage, key ID, val int)

@[c: 'ImGuiStorage_GetBool']
fn storage_get_bool(self &Storage, key ID, default_val bool) bool

@[c: 'ImGuiStorage_SetBool']
fn storage_set_bool(self &Storage, key ID, val bool)

@[c: 'ImGuiStorage_GetFloat']
fn storage_get_float(self &Storage, key ID, default_val f32) f32

@[c: 'ImGuiStorage_SetFloat']
fn storage_set_float(self &Storage, key ID, val f32)

@[c: 'ImGuiStorage_GetVoidPtr']
fn storage_get_void_ptr(self &Storage, key ID) voidptr

@[c: 'ImGuiStorage_SetVoidPtr']
fn storage_set_void_ptr(self &Storage, key ID, val voidptr)

@[c: 'ImGuiStorage_GetIntRef']
fn storage_get_int_ref(self &Storage, key ID, default_val int) &int

@[c: 'ImGuiStorage_GetBoolRef']
fn storage_get_bool_ref(self &Storage, key ID, default_val bool) &bool

@[c: 'ImGuiStorage_GetFloatRef']
fn storage_get_float_ref(self &Storage, key ID, default_val f32) &f32

@[c: 'ImGuiStorage_GetVoidPtrRef']
fn storage_get_void_ptr_ref(self &Storage, key ID, default_val voidptr) &voidptr

@[c: 'ImGuiStorage_BuildSortByKey']
fn storage_build_sort_by_key(self &Storage)

@[c: 'ImGuiStorage_SetAllInt']
fn storage_set_all_int(self &Storage, val int)

@[c: 'ImGuiListClipper_ImGuiListClipper']
fn list_clipper_im_gui_list_clipper() &ListClipper

@[c: 'ImGuiListClipper_ImGuiListClipper_Construct']
fn list_clipper_im_gui_list_clipper_construct(self &ListClipper)

@[c: 'ImGuiListClipper_destroy']
fn list_clipper_destroy(self &ListClipper)

@[c: 'ImGuiListClipper_Begin']
fn list_clipper_begin(self &ListClipper, items_count int, items_height f32)

@[c: 'ImGuiListClipper_End']
fn list_clipper_end(self &ListClipper)

@[c: 'ImGuiListClipper_Step']
fn list_clipper_step(self &ListClipper) bool

@[c: 'ImGuiListClipper_IncludeItemByIndex']
fn list_clipper_include_item_by_index(self &ListClipper, item_index int)

@[c: 'ImGuiListClipper_IncludeItemsByIndex']
fn list_clipper_include_items_by_index(self &ListClipper, item_begin int, item_end int)

@[c: 'ImGuiListClipper_SeekCursorForItem']
fn list_clipper_seek_cursor_for_item(self &ListClipper, item_index int)

@[c: 'ImColor_ImColor_Nil']
fn im_color_im_color_nil() &ImColor

@[c: 'ImColor_ImColor_Nil_Construct']
fn im_color_im_color_nil_construct(self &ImColor)

@[c: 'ImColor_destroy']
fn im_color_destroy(self &ImColor)

@[c: 'ImColor_ImColor_Float']
fn im_color_im_color_float(r f32, g f32, b f32, a f32) &ImColor

@[c: 'ImColor_ImColor_Float_Construct']
fn im_color_im_color_float_construct(self &ImColor, r f32, g f32, b f32, a f32)

@[c: 'ImColor_ImColor_Vec4']
fn im_color_im_color_vec4(col C.ImVec4) &ImColor

@[c: 'ImColor_ImColor_Vec4_Construct']
fn im_color_im_color_vec4_construct(self &ImColor, col C.ImVec4)

@[c: 'ImColor_ImColor_Int']
fn im_color_im_color_int(r int, g int, b int, a int) &ImColor

@[c: 'ImColor_ImColor_Int_Construct']
fn im_color_im_color_int_construct(self &ImColor, r int, g int, b int, a int)

@[c: 'ImColor_ImColor_U32']
fn im_color_im_color_u32(rgba ImU32) &ImColor

@[c: 'ImColor_ImColor_U32_Construct']
fn im_color_im_color_u32_construct(self &ImColor, rgba ImU32)

@[c: 'ImColor_SetHSV']
fn im_color_set_hsv(self &ImColor, h f32, s f32, v f32, a f32)

@[c: 'ImColor_HSV']
fn im_color_hsv(p_out &ImColor, h f32, s f32, v f32, a f32)

@[c: 'ImGuiSelectionBasicStorage_ImGuiSelectionBasicStorage']
fn selection_basic_storage_im_gui_selection_basic_storage() &SelectionBasicStorage

@[c: 'ImGuiSelectionBasicStorage_ImGuiSelectionBasicStorage_Construct']
fn selection_basic_storage_im_gui_selection_basic_storage_construct(self &SelectionBasicStorage)

@[c: 'ImGuiSelectionBasicStorage_destroy']
fn selection_basic_storage_destroy(self &SelectionBasicStorage)

@[c: 'ImGuiSelectionBasicStorage_ApplyRequests']
fn selection_basic_storage_apply_requests(self &SelectionBasicStorage, ms_io &MultiSelectIO)

@[c: 'ImGuiSelectionBasicStorage_Contains']
fn selection_basic_storage_contains(self &SelectionBasicStorage, id ID) bool

@[c: 'ImGuiSelectionBasicStorage_Clear']
fn selection_basic_storage_clear(self &SelectionBasicStorage)

@[c: 'ImGuiSelectionBasicStorage_Swap']
fn selection_basic_storage_swap(self &SelectionBasicStorage, r &SelectionBasicStorage)

@[c: 'ImGuiSelectionBasicStorage_SetItemSelected']
fn selection_basic_storage_set_item_selected(self &SelectionBasicStorage, id ID, selected bool)

@[c: 'ImGuiSelectionBasicStorage_GetNextSelectedItem']
fn selection_basic_storage_get_next_selected_item(self &SelectionBasicStorage, opaque_it &voidptr, out_id &ID) bool

@[c: 'ImGuiSelectionBasicStorage_GetStorageIdFromIndex']
fn selection_basic_storage_get_storage_id_from_index(self &SelectionBasicStorage, idx int) ID

@[c: 'ImGuiSelectionExternalStorage_ImGuiSelectionExternalStorage']
fn selection_external_storage_im_gui_selection_external_storage() &C.ImGuiSelectionExternalStorage

@[c: 'ImGuiSelectionExternalStorage_ImGuiSelectionExternalStorage_Construct']
fn selection_external_storage_im_gui_selection_external_storage_construct(self &C.ImGuiSelectionExternalStorage)

@[c: 'ImGuiSelectionExternalStorage_destroy']
fn selection_external_storage_destroy(self &C.ImGuiSelectionExternalStorage)

@[c: 'ImGuiSelectionExternalStorage_ApplyRequests']
fn selection_external_storage_apply_requests(self &C.ImGuiSelectionExternalStorage, ms_io &MultiSelectIO)

@[c: 'ImDrawCmd_ImDrawCmd']
fn im_draw_cmd_im_draw_cmd() &ImDrawCmd

@[c: 'ImDrawCmd_ImDrawCmd_Construct']
fn im_draw_cmd_im_draw_cmd_construct(self &ImDrawCmd)

@[c: 'ImDrawCmd_destroy']
fn im_draw_cmd_destroy(self &ImDrawCmd)

@[c: 'ImDrawCmd_GetTexID']
fn im_draw_cmd_get_tex_id(self &ImDrawCmd) ImTextureID

@[c: 'ImDrawListSplitter_ImDrawListSplitter']
fn im_draw_list_splitter_im_draw_list_splitter() &ImDrawListSplitter

@[c: 'ImDrawListSplitter_ImDrawListSplitter_Construct']
fn im_draw_list_splitter_im_draw_list_splitter_construct(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_destroy']
fn im_draw_list_splitter_destroy(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_Clear']
fn im_draw_list_splitter_clear(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_ClearFreeMemory']
fn im_draw_list_splitter_clear_free_memory(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_Split']
fn im_draw_list_splitter_split(self &ImDrawListSplitter, draw_list &ImDrawList, count int)

@[c: 'ImDrawListSplitter_Merge']
fn im_draw_list_splitter_merge(self &ImDrawListSplitter, draw_list &ImDrawList)

@[c: 'ImDrawListSplitter_SetCurrentChannel']
fn im_draw_list_splitter_set_current_channel(self &ImDrawListSplitter, draw_list &ImDrawList, channel_idx int)

@[c: 'ImDrawList_ImDrawList']
fn im_draw_list_im_draw_list(shared_data &ImDrawListSharedData) &ImDrawList

@[c: 'ImDrawList_ImDrawList_Construct']
fn im_draw_list_im_draw_list_construct(self &ImDrawList, shared_data &ImDrawListSharedData)

@[c: 'ImDrawList_destroy']
fn im_draw_list_destroy(self &ImDrawList)

@[c: 'ImDrawList_PushClipRect']
fn im_draw_list_push_clip_rect(self &ImDrawList, clip_rect_min ImVec2, clip_rect_max ImVec2, intersect_with_current_clip_rect bool)

@[c: 'ImDrawList_PushClipRectFullScreen']
fn im_draw_list_push_clip_rect_full_screen(self &ImDrawList)

@[c: 'ImDrawList_PopClipRect']
fn im_draw_list_pop_clip_rect(self &ImDrawList)

@[c: 'ImDrawList_PushTextureID']
fn im_draw_list_push_texture_id(self &ImDrawList, texture_id ImTextureID)

@[c: 'ImDrawList_PopTextureID']
fn im_draw_list_pop_texture_id(self &ImDrawList)

@[c: 'ImDrawList_GetClipRectMin']
fn im_draw_list_get_clip_rect_min(p_out &ImVec2, self &ImDrawList)

@[c: 'ImDrawList_GetClipRectMax']
fn im_draw_list_get_clip_rect_max(p_out &ImVec2, self &ImDrawList)

@[c: 'ImDrawList_AddLine']
fn im_draw_list_add_line(self &ImDrawList, p1 ImVec2, p2 ImVec2, col ImU32, thickness f32)

@[c: 'ImDrawList_AddRect']
fn im_draw_list_add_rect(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags, thickness f32)

@[c: 'ImDrawList_AddRectFilled']
fn im_draw_list_add_rect_filled(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags)

@[c: 'ImDrawList_AddRectFilledMultiColor']
fn im_draw_list_add_rect_filled_multi_color(self &ImDrawList, p_min ImVec2, p_max ImVec2, col_upr_left ImU32, col_upr_right ImU32, col_bot_right ImU32, col_bot_left ImU32)

@[c: 'ImDrawList_AddQuad']
fn im_draw_list_add_quad(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32, thickness f32)

@[c: 'ImDrawList_AddQuadFilled']
fn im_draw_list_add_quad_filled(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32)

@[c: 'ImDrawList_AddTriangle']
fn im_draw_list_add_triangle(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32, thickness f32)

@[c: 'ImDrawList_AddTriangleFilled']
fn im_draw_list_add_triangle_filled(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32)

@[c: 'ImDrawList_AddCircle']
fn im_draw_list_add_circle(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int, thickness f32)

@[c: 'ImDrawList_AddCircleFilled']
fn im_draw_list_add_circle_filled(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

@[c: 'ImDrawList_AddNgon']
fn im_draw_list_add_ngon(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int, thickness f32)

@[c: 'ImDrawList_AddNgonFilled']
fn im_draw_list_add_ngon_filled(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

@[c: 'ImDrawList_AddEllipse']
fn im_draw_list_add_ellipse(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32, rot f32, num_segments int, thickness f32)

@[c: 'ImDrawList_AddEllipseFilled']
fn im_draw_list_add_ellipse_filled(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32, rot f32, num_segments int)

@[c: 'ImDrawList_AddText_Vec2']
fn im_draw_list_add_text_vec2(self &ImDrawList, pos ImVec2, col ImU32, text_begin &i8, text_end &i8)

@[c: 'ImDrawList_AddText_FontPtr']
fn im_draw_list_add_text_font_ptr(self &ImDrawList, font &ImFont, font_size f32, pos ImVec2, col ImU32, text_begin &i8, text_end &i8, wrap_width f32, cpu_fine_clip_rect &C.ImVec4)

@[c: 'ImDrawList_AddBezierCubic']
fn im_draw_list_add_bezier_cubic(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32, thickness f32, num_segments int)

@[c: 'ImDrawList_AddBezierQuadratic']
fn im_draw_list_add_bezier_quadratic(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32, thickness f32, num_segments int)

@[c: 'ImDrawList_AddPolyline']
fn im_draw_list_add_polyline(self &ImDrawList, points &ImVec2, num_points int, col ImU32, flags ImDrawFlags, thickness f32)

@[c: 'ImDrawList_AddConvexPolyFilled']
fn im_draw_list_add_convex_poly_filled(self &ImDrawList, points &ImVec2, num_points int, col ImU32)

@[c: 'ImDrawList_AddConcavePolyFilled']
fn im_draw_list_add_concave_poly_filled(self &ImDrawList, points &ImVec2, num_points int, col ImU32)

@[c: 'ImDrawList_AddImage']
fn im_draw_list_add_image(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2, uv_min ImVec2, uv_max ImVec2, col ImU32)

@[c: 'ImDrawList_AddImageQuad']
fn im_draw_list_add_image_quad(self &ImDrawList, user_texture_id ImTextureID, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, uv1 ImVec2, uv2 ImVec2, uv3 ImVec2, uv4 ImVec2, col ImU32)

@[c: 'ImDrawList_AddImageRounded']
fn im_draw_list_add_image_rounded(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2, uv_min ImVec2, uv_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags)

@[c: 'ImDrawList_PathClear']
fn im_draw_list_path_clear(self &ImDrawList)

@[c: 'ImDrawList_PathLineTo']
fn im_draw_list_path_line_to(self &ImDrawList, pos ImVec2)

@[c: 'ImDrawList_PathLineToMergeDuplicate']
fn im_draw_list_path_line_to_merge_duplicate(self &ImDrawList, pos ImVec2)

@[c: 'ImDrawList_PathFillConvex']
fn im_draw_list_path_fill_convex(self &ImDrawList, col ImU32)

@[c: 'ImDrawList_PathFillConcave']
fn im_draw_list_path_fill_concave(self &ImDrawList, col ImU32)

@[c: 'ImDrawList_PathStroke']
fn im_draw_list_path_stroke(self &ImDrawList, col ImU32, flags ImDrawFlags, thickness f32)

@[c: 'ImDrawList_PathArcTo']
fn im_draw_list_path_arc_to(self &ImDrawList, center ImVec2, radius f32, a_min f32, a_max f32, num_segments int)

@[c: 'ImDrawList_PathArcToFast']
fn im_draw_list_path_arc_to_fast(self &ImDrawList, center ImVec2, radius f32, a_min_of_12 int, a_max_of_12 int)

@[c: 'ImDrawList_PathEllipticalArcTo']
fn im_draw_list_path_elliptical_arc_to(self &ImDrawList, center ImVec2, radius ImVec2, rot f32, a_min f32, a_max f32, num_segments int)

@[c: 'ImDrawList_PathBezierCubicCurveTo']
fn im_draw_list_path_bezier_cubic_curve_to(self &ImDrawList, p2 ImVec2, p3 ImVec2, p4 ImVec2, num_segments int)

@[c: 'ImDrawList_PathBezierQuadraticCurveTo']
fn im_draw_list_path_bezier_quadratic_curve_to(self &ImDrawList, p2 ImVec2, p3 ImVec2, num_segments int)

@[c: 'ImDrawList_PathRect']
fn im_draw_list_path_rect(self &ImDrawList, rect_min ImVec2, rect_max ImVec2, rounding f32, flags ImDrawFlags)

@[c: 'ImDrawList_AddCallback']
fn im_draw_list_add_callback(self &ImDrawList, callback ImDrawCallback, userdata voidptr, userdata_size usize)

@[c: 'ImDrawList_AddDrawCmd']
fn im_draw_list_add_draw_cmd(self &ImDrawList)

@[c: 'ImDrawList_CloneOutput']
fn im_draw_list_clone_output(self &ImDrawList) &ImDrawList

@[c: 'ImDrawList_ChannelsSplit']
fn im_draw_list_channels_split(self &ImDrawList, count int)

@[c: 'ImDrawList_ChannelsMerge']
fn im_draw_list_channels_merge(self &ImDrawList)

@[c: 'ImDrawList_ChannelsSetCurrent']
fn im_draw_list_channels_set_current(self &ImDrawList, n int)

@[c: 'ImDrawList_PrimReserve']
fn im_draw_list_prim_reserve(self &ImDrawList, idx_count int, vtx_count int)

@[c: 'ImDrawList_PrimUnreserve']
fn im_draw_list_prim_unreserve(self &ImDrawList, idx_count int, vtx_count int)

@[c: 'ImDrawList_PrimRect']
fn im_draw_list_prim_rect(self &ImDrawList, a ImVec2, b ImVec2, col ImU32)

@[c: 'ImDrawList_PrimRectUV']
fn im_draw_list_prim_rect_uv(self &ImDrawList, a ImVec2, b ImVec2, uv_a ImVec2, uv_b ImVec2, col ImU32)

@[c: 'ImDrawList_PrimQuadUV']
fn im_draw_list_prim_quad_uv(self &ImDrawList, a ImVec2, b ImVec2, c ImVec2, d ImVec2, uv_a ImVec2, uv_b ImVec2, uv_c ImVec2, uv_d ImVec2, col ImU32)

@[c: 'ImDrawList_PrimWriteVtx']
fn im_draw_list_prim_write_vtx(self &ImDrawList, pos ImVec2, uv ImVec2, col ImU32)

@[c: 'ImDrawList_PrimWriteIdx']
fn im_draw_list_prim_write_idx(self &ImDrawList, idx ImDrawIdx)

@[c: 'ImDrawList_PrimVtx']
fn im_draw_list_prim_vtx(self &ImDrawList, pos ImVec2, uv ImVec2, col ImU32)

@[c: 'ImDrawList__ResetForNewFrame']
fn im_draw_list__reset_for_new_frame(self &ImDrawList)

@[c: 'ImDrawList__ClearFreeMemory']
fn im_draw_list__clear_free_memory(self &ImDrawList)

@[c: 'ImDrawList__PopUnusedDrawCmd']
fn im_draw_list__pop_unused_draw_cmd(self &ImDrawList)

@[c: 'ImDrawList__TryMergeDrawCmds']
fn im_draw_list__try_merge_draw_cmds(self &ImDrawList)

@[c: 'ImDrawList__OnChangedClipRect']
fn im_draw_list__on_changed_clip_rect(self &ImDrawList)

@[c: 'ImDrawList__OnChangedTextureID']
fn im_draw_list__on_changed_texture_id(self &ImDrawList)

@[c: 'ImDrawList__OnChangedVtxOffset']
fn im_draw_list__on_changed_vtx_offset(self &ImDrawList)

@[c: 'ImDrawList__SetTextureID']
fn im_draw_list__set_texture_id(self &ImDrawList, texture_id ImTextureID)

@[c: 'ImDrawList__CalcCircleAutoSegmentCount']
fn im_draw_list__calc_circle_auto_segment_count(self &ImDrawList, radius f32) int

@[c: 'ImDrawList__PathArcToFastEx']
fn im_draw_list__path_arc_to_fast_ex(self &ImDrawList, center ImVec2, radius f32, a_min_sample int, a_max_sample int, a_step int)

@[c: 'ImDrawList__PathArcToN']
fn im_draw_list__path_arc_to_n(self &ImDrawList, center ImVec2, radius f32, a_min f32, a_max f32, num_segments int)

@[c: 'ImDrawData_ImDrawData']
fn im_draw_data_im_draw_data() &ImDrawData

@[c: 'ImDrawData_ImDrawData_Construct']
fn im_draw_data_im_draw_data_construct(self &ImDrawData)

@[c: 'ImDrawData_destroy']
fn im_draw_data_destroy(self &ImDrawData)

@[c: 'ImDrawData_Clear']
fn im_draw_data_clear(self &ImDrawData)

@[c: 'ImDrawData_AddDrawList']
fn im_draw_data_add_draw_list(self &ImDrawData, draw_list &ImDrawList)

@[c: 'ImDrawData_DeIndexAllBuffers']
fn im_draw_data_de_index_all_buffers(self &ImDrawData)

@[c: 'ImDrawData_ScaleClipRects']
fn im_draw_data_scale_clip_rects(self &ImDrawData, fb_scale ImVec2)

@[c: 'ImFontConfig_ImFontConfig']
fn im_font_config_im_font_config() &ImFontConfig

@[c: 'ImFontConfig_ImFontConfig_Construct']
fn im_font_config_im_font_config_construct(self &ImFontConfig)

@[c: 'ImFontConfig_destroy']
fn im_font_config_destroy(self &ImFontConfig)

@[c: 'ImFontGlyphRangesBuilder_ImFontGlyphRangesBuilder']
fn im_font_glyph_ranges_builder_im_font_glyph_ranges_builder() &ImFontGlyphRangesBuilder

@[c: 'ImFontGlyphRangesBuilder_ImFontGlyphRangesBuilder_Construct']
fn im_font_glyph_ranges_builder_im_font_glyph_ranges_builder_construct(self &ImFontGlyphRangesBuilder)

@[c: 'ImFontGlyphRangesBuilder_destroy']
fn im_font_glyph_ranges_builder_destroy(self &ImFontGlyphRangesBuilder)

@[c: 'ImFontGlyphRangesBuilder_Clear']
fn im_font_glyph_ranges_builder_clear(self &ImFontGlyphRangesBuilder)

@[c: 'ImFontGlyphRangesBuilder_GetBit']
fn im_font_glyph_ranges_builder_get_bit(self &ImFontGlyphRangesBuilder, n usize) bool

@[c: 'ImFontGlyphRangesBuilder_SetBit']
fn im_font_glyph_ranges_builder_set_bit(self &ImFontGlyphRangesBuilder, n usize)

@[c: 'ImFontGlyphRangesBuilder_AddChar']
fn im_font_glyph_ranges_builder_add_char(self &ImFontGlyphRangesBuilder, c C.ImWchar)

@[c: 'ImFontGlyphRangesBuilder_AddText']
fn im_font_glyph_ranges_builder_add_text(self &ImFontGlyphRangesBuilder, text &i8, text_end &i8)

@[c: 'ImFontGlyphRangesBuilder_AddRanges']
fn im_font_glyph_ranges_builder_add_ranges(self &ImFontGlyphRangesBuilder, ranges &C.ImWchar)

@[c: 'ImFontGlyphRangesBuilder_BuildRanges']
fn im_font_glyph_ranges_builder_build_ranges(self &ImFontGlyphRangesBuilder, out_ranges &ImVector_ImWchar)

@[c: 'ImFontAtlasCustomRect_ImFontAtlasCustomRect']
fn im_font_atlas_custom_rect_im_font_atlas_custom_rect() &ImFontAtlasCustomRect

@[c: 'ImFontAtlasCustomRect_ImFontAtlasCustomRect_Construct']
fn im_font_atlas_custom_rect_im_font_atlas_custom_rect_construct(self &ImFontAtlasCustomRect)

@[c: 'ImFontAtlasCustomRect_destroy']
fn im_font_atlas_custom_rect_destroy(self &ImFontAtlasCustomRect)

@[c: 'ImFontAtlasCustomRect_IsPacked']
fn im_font_atlas_custom_rect_is_packed(self &ImFontAtlasCustomRect) bool

@[c: 'ImFontAtlas_ImFontAtlas']
fn im_font_atlas_im_font_atlas() &ImFontAtlas

@[c: 'ImFontAtlas_ImFontAtlas_Construct']
fn im_font_atlas_im_font_atlas_construct(self &ImFontAtlas)

@[c: 'ImFontAtlas_destroy']
fn im_font_atlas_destroy(self &ImFontAtlas)

@[c: 'ImFontAtlas_AddFont']
fn im_font_atlas_add_font(self &ImFontAtlas, font_cfg &ImFontConfig) &ImFont

@[c: 'ImFontAtlas_AddFontDefault']
fn im_font_atlas_add_font_default(self &ImFontAtlas, font_cfg &ImFontConfig) &ImFont

@[c: 'ImFontAtlas_AddFontFromFileTTF']
fn im_font_atlas_add_font_from_file_ttf(self &ImFontAtlas, filename &i8, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

@[c: 'ImFontAtlas_AddFontFromMemoryTTF']
fn im_font_atlas_add_font_from_memory_ttf(self &ImFontAtlas, font_data voidptr, font_data_size int, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

@[c: 'ImFontAtlas_AddFontFromMemoryCompressedTTF']
fn im_font_atlas_add_font_from_memory_compressed_ttf(self &ImFontAtlas, compressed_font_data voidptr, compressed_font_data_size int, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

@[c: 'ImFontAtlas_AddFontFromMemoryCompressedBase85TTF']
fn im_font_atlas_add_font_from_memory_compressed_base85_ttf(self &ImFontAtlas, compressed_font_data_base85 &i8, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

@[c: 'ImFontAtlas_ClearInputData']
fn im_font_atlas_clear_input_data(self &ImFontAtlas)

@[c: 'ImFontAtlas_ClearFonts']
fn im_font_atlas_clear_fonts(self &ImFontAtlas)

@[c: 'ImFontAtlas_ClearTexData']
fn im_font_atlas_clear_tex_data(self &ImFontAtlas)

@[c: 'ImFontAtlas_Clear']
fn im_font_atlas_clear(self &ImFontAtlas)

@[c: 'ImFontAtlas_Build']
fn im_font_atlas_build(self &ImFontAtlas) bool

@[c: 'ImFontAtlas_GetTexDataAsAlpha8']
fn im_font_atlas_get_tex_data_as_alpha8(self &ImFontAtlas, out_pixels &&u8, out_width &int, out_height &int, out_bytes_per_pixel &int)

@[c: 'ImFontAtlas_GetTexDataAsRGBA32']
fn im_font_atlas_get_tex_data_as_rgba_32(self &ImFontAtlas, out_pixels &&u8, out_width &int, out_height &int, out_bytes_per_pixel &int)

@[c: 'ImFontAtlas_IsBuilt']
fn im_font_atlas_is_built(self &ImFontAtlas) bool

@[c: 'ImFontAtlas_SetTexID']
fn im_font_atlas_set_tex_id(self &ImFontAtlas, id ImTextureID)

@[c: 'ImFontAtlas_GetGlyphRangesDefault']
fn im_font_atlas_get_glyph_ranges_default(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesGreek']
fn im_font_atlas_get_glyph_ranges_greek(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesKorean']
fn im_font_atlas_get_glyph_ranges_korean(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesJapanese']
fn im_font_atlas_get_glyph_ranges_japanese(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesChineseFull']
fn im_font_atlas_get_glyph_ranges_chinese_full(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesChineseSimplifiedCommon']
fn im_font_atlas_get_glyph_ranges_chinese_simplified_common(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesCyrillic']
fn im_font_atlas_get_glyph_ranges_cyrillic(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesThai']
fn im_font_atlas_get_glyph_ranges_thai(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesVietnamese']
fn im_font_atlas_get_glyph_ranges_vietnamese(self &ImFontAtlas) &C.ImWchar

@[c: 'ImFontAtlas_AddCustomRectRegular']
fn im_font_atlas_add_custom_rect_regular(self &ImFontAtlas, width int, height int) int

@[c: 'ImFontAtlas_AddCustomRectFontGlyph']
fn im_font_atlas_add_custom_rect_font_glyph(self &ImFontAtlas, font &ImFont, id C.ImWchar, width int, height int, advance_x f32, offset ImVec2) int

@[c: 'ImFontAtlas_GetCustomRectByIndex']
fn im_font_atlas_get_custom_rect_by_index(self &ImFontAtlas, index int) &ImFontAtlasCustomRect

@[c: 'ImFontAtlas_CalcCustomRectUV']
fn im_font_atlas_calc_custom_rect_uv(self &ImFontAtlas, rect &ImFontAtlasCustomRect, out_uv_min &ImVec2, out_uv_max &ImVec2)

@[c: 'ImFont_ImFont']
fn im_font_im_font() &ImFont

@[c: 'ImFont_ImFont_Construct']
fn im_font_im_font_construct(self &ImFont)

@[c: 'ImFont_destroy']
fn im_font_destroy(self &ImFont)

@[c: 'ImFont_FindGlyph']
fn im_font_find_glyph(self &ImFont, c C.ImWchar) &ImFontGlyph

@[c: 'ImFont_FindGlyphNoFallback']
fn im_font_find_glyph_no_fallback(self &ImFont, c C.ImWchar) &ImFontGlyph

@[c: 'ImFont_GetCharAdvance']
fn im_font_get_char_advance(self &ImFont, c C.ImWchar) f32

@[c: 'ImFont_IsLoaded']
fn im_font_is_loaded(self &ImFont) bool

@[c: 'ImFont_GetDebugName']
fn im_font_get_debug_name(self &ImFont) &i8

@[c: 'ImFont_CalcTextSizeA']
fn im_font_calc_text_size_a(p_out &ImVec2, self &ImFont, size f32, max_width f32, wrap_width f32, text_begin &i8, text_end &i8, remaining &&u8)

@[c: 'ImFont_CalcWordWrapPositionA']
fn im_font_calc_word_wrap_position_a(self &ImFont, scale f32, text &i8, text_end &i8, wrap_width f32) &i8

@[c: 'ImFont_RenderChar']
fn im_font_render_char(self &ImFont, draw_list &ImDrawList, size f32, pos ImVec2, col ImU32, c C.ImWchar)

@[c: 'ImFont_RenderText']
fn im_font_render_text(self &ImFont, draw_list &ImDrawList, size f32, pos ImVec2, col ImU32, clip_rect C.ImVec4, text_begin &i8, text_end &i8, wrap_width f32, cpu_fine_clip bool)

@[c: 'ImFont_BuildLookupTable']
fn im_font_build_lookup_table(self &ImFont)

@[c: 'ImFont_ClearOutputData']
fn im_font_clear_output_data(self &ImFont)

@[c: 'ImFont_GrowIndex']
fn im_font_grow_index(self &ImFont, new_size int)

@[c: 'ImFont_AddGlyph']
fn im_font_add_glyph(self &ImFont, src_cfg &ImFontConfig, c C.ImWchar, x0 f32, y0 f32, x1 f32, y1 f32, u0 f32, v0 f32, u1 f32, v1 f32, advance_x f32)

@[c: 'ImFont_AddRemapChar']
fn im_font_add_remap_char(self &ImFont, dst C.ImWchar, src C.ImWchar, overwrite_dst bool)

@[c: 'ImFont_IsGlyphRangeUnused']
fn im_font_is_glyph_range_unused(self &ImFont, c_begin u32, c_last u32) bool

@[c: 'ImGuiViewport_ImGuiViewport']
fn viewport_im_gui_viewport() &Viewport

@[c: 'ImGuiViewport_ImGuiViewport_Construct']
fn viewport_im_gui_viewport_construct(self &Viewport)

@[c: 'ImGuiViewport_destroy']
fn viewport_destroy(self &Viewport)

@[c: 'ImGuiViewport_GetCenter']
fn viewport_get_center(p_out &ImVec2, self &Viewport)

@[c: 'ImGuiViewport_GetWorkCenter']
fn viewport_get_work_center(p_out &ImVec2, self &Viewport)

@[c: 'ImGuiPlatformIO_ImGuiPlatformIO']
fn platform_io_im_gui_platform_io() &PlatformIO

@[c: 'ImGuiPlatformIO_ImGuiPlatformIO_Construct']
fn platform_io_im_gui_platform_io_construct(self &PlatformIO)

@[c: 'ImGuiPlatformIO_destroy']
fn platform_io_destroy(self &PlatformIO)

@[c: 'ImGuiPlatformMonitor_ImGuiPlatformMonitor']
fn platform_monitor_im_gui_platform_monitor() &PlatformMonitor

@[c: 'ImGuiPlatformMonitor_ImGuiPlatformMonitor_Construct']
fn platform_monitor_im_gui_platform_monitor_construct(self &PlatformMonitor)

@[c: 'ImGuiPlatformMonitor_destroy']
fn platform_monitor_destroy(self &PlatformMonitor)

@[c: 'ImGuiPlatformImeData_ImGuiPlatformImeData']
fn platform_ime_data_im_gui_platform_ime_data() &PlatformImeData

@[c: 'ImGuiPlatformImeData_ImGuiPlatformImeData_Construct']
fn platform_ime_data_im_gui_platform_ime_data_construct(self &PlatformImeData)

@[c: 'ImGuiPlatformImeData_destroy']
fn platform_ime_data_destroy(self &PlatformImeData)

@[c: 'igImHashData']
fn im_hash_data(data voidptr, data_size usize, seed ID) ID

@[c: 'igImHashStr']
fn im_hash_str(data &i8, data_size usize, seed ID) ID

@[c: 'igImQsort']
fn im_qsort(base voidptr, count usize, size_of_element usize, compare_func fn (voidptr, voidptr) int)

@[c: 'igImAlphaBlendColors']
fn im_alpha_blend_colors(col_a ImU32, col_b ImU32) ImU32

@[c: 'igImIsPowerOfTwo_Int']
fn im_is_power_of_two_int(v int) bool

@[c: 'igImIsPowerOfTwo_U64']
fn im_is_power_of_two_u64(v ImU64) bool

@[c: 'igImUpperPowerOfTwo']
fn im_upper_power_of_two(v int) int

@[c: 'igImCountSetBits']
fn im_count_set_bits(v u32) u32

@[c: 'igImStricmp']
fn im_stricmp(str1 &i8, str2 &i8) int

@[c: 'igImStrnicmp']
fn im_strnicmp(str1 &i8, str2 &i8, count usize) int

@[c: 'igImStrncpy']
fn im_strncpy(dst &i8, src &i8, count usize)

@[c: 'igImStrdup']
fn im_strdup(str &i8) &i8

@[c: 'igImStrdupcpy']
fn im_strdupcpy(dst &i8, p_dst_size &usize, str &i8) &i8

@[c: 'igImStrchrRange']
fn im_strchr_range(str_begin &i8, str_end &i8, c i8) &i8

@[c: 'igImStreolRange']
fn im_streol_range(str &i8, str_end &i8) &i8

@[c: 'igImStristr']
fn im_stristr(haystack &i8, haystack_end &i8, needle &i8, needle_end &i8) &i8

@[c: 'igImStrTrimBlanks']
fn im_str_trim_blanks(str &i8)

@[c: 'igImStrSkipBlank']
fn im_str_skip_blank(str &i8) &i8

@[c: 'igImStrlenW']
fn im_strlen_w(str &C.ImWchar) int

@[c: 'igImStrbol']
fn im_strbol(buf_mid_line &i8, buf_begin &i8) &i8

@[c: 'igImToUpper']
fn im_to_upper(c i8) i8

@[c: 'igImCharIsBlankA']
fn im_char_is_blank_a(c i8) bool

@[c: 'igImCharIsBlankW']
fn im_char_is_blank_w(c u32) bool

@[c: 'igImCharIsXdigitA']
fn im_char_is_xdigit_a(c i8) bool

@[c: 'igImFormatString']
@[c2v_variadic]
fn im_format_string(buf &i8, buf_size usize, fmt ...&i8) int

@[c: 'igImFormatStringV']
fn im_format_string_v(buf &i8, buf_size usize, fmt &i8, args C.va_list) int

@[c: 'igImFormatStringToTempBuffer']
@[c2v_variadic]
fn im_format_string_to_temp_buffer(out_buf &&u8, out_buf_end &&u8, fmt ...&i8)

@[c: 'igImFormatStringToTempBufferV']
fn im_format_string_to_temp_buffer_v(out_buf &&u8, out_buf_end &&u8, fmt &i8, args C.va_list)

@[c: 'igImParseFormatFindStart']
fn im_parse_format_find_start(format &i8) &i8

@[c: 'igImParseFormatFindEnd']
fn im_parse_format_find_end(format &i8) &i8

@[c: 'igImParseFormatTrimDecorations']
fn im_parse_format_trim_decorations(format &i8, buf &i8, buf_size usize) &i8

@[c: 'igImParseFormatSanitizeForPrinting']
fn im_parse_format_sanitize_for_printing(fmt_in &i8, fmt_out &i8, fmt_out_size usize)

@[c: 'igImParseFormatSanitizeForScanning']
fn im_parse_format_sanitize_for_scanning(fmt_in &i8, fmt_out &i8, fmt_out_size usize) &i8

@[c: 'igImParseFormatPrecision']
fn im_parse_format_precision(format &i8, default_value int) int

@[c: 'igImTextCharToUtf8']
fn im_text_char_to_utf8(out_buf &i8, c u32) &i8

@[c: 'igImTextStrToUtf8']
fn im_text_str_to_utf8(out_buf &i8, out_buf_size int, in_text &C.ImWchar, in_text_end &C.ImWchar) int

@[c: 'igImTextCharFromUtf8']
fn im_text_char_from_utf8(out_char &u32, in_text &i8, in_text_end &i8) int

@[c: 'igImTextStrFromUtf8']
fn im_text_str_from_utf8(out_buf &C.ImWchar, out_buf_size int, in_text &i8, in_text_end &i8, in_remaining &&u8) int

@[c: 'igImTextCountCharsFromUtf8']
fn im_text_count_chars_from_utf8(in_text &i8, in_text_end &i8) int

@[c: 'igImTextCountUtf8BytesFromChar']
fn im_text_count_utf8_bytes_from_char(in_text &i8, in_text_end &i8) int

@[c: 'igImTextCountUtf8BytesFromStr']
fn im_text_count_utf8_bytes_from_str(in_text &C.ImWchar, in_text_end &C.ImWchar) int

@[c: 'igImTextFindPreviousUtf8Codepoint']
fn im_text_find_previous_utf8_codepoint(in_text_start &i8, in_text_curr &i8) &i8

@[c: 'igImTextCountLines']
fn im_text_count_lines(in_text &i8, in_text_end &i8) int

@[c: 'igImFileOpen']
fn im_file_open(filename &i8, mode &i8) ImFileHandle

@[c: 'igImFileClose']
fn im_file_close(file ImFileHandle) bool

@[c: 'igImFileGetSize']
fn im_file_get_size(file ImFileHandle) ImU64

@[c: 'igImFileRead']
fn im_file_read(data voidptr, size ImU64, count ImU64, file ImFileHandle) ImU64

@[c: 'igImFileWrite']
fn im_file_write(data voidptr, size ImU64, count ImU64, file ImFileHandle) ImU64

@[c: 'igImFileLoadToMemory']
fn im_file_load_to_memory(filename &i8, mode &i8, out_file_size &usize, padding_bytes int) voidptr

@[c: 'igImPow_Float']
fn im_pow_float(x f32, y f32) f32

@[c: 'igImPow_double']
fn im_pow_double(x f64, y f64) f64

@[c: 'igImLog_Float']
fn im_log_float(x f32) f32

@[c: 'igImLog_double']
fn im_log_double(x f64) f64

@[c: 'igImAbs_Int']
fn im_abs_int(x int) int

@[c: 'igImAbs_Float']
fn im_abs_float(x f32) f32

@[c: 'igImAbs_double']
fn im_abs_double(x f64) f64

@[c: 'igImSign_Float']
fn im_sign_float(x f32) f32

@[c: 'igImSign_double']
fn im_sign_double(x f64) f64

@[c: 'igImRsqrt_Float']
fn im_rsqrt_float(x f32) f32

@[c: 'igImRsqrt_double']
fn im_rsqrt_double(x f64) f64

@[c: 'igImMin']
fn im_min(p_out &ImVec2, lhs ImVec2, rhs ImVec2)

@[c: 'igImMax']
fn im_max(p_out &ImVec2, lhs ImVec2, rhs ImVec2)

@[c: 'igImClamp']
fn im_clamp(p_out &ImVec2, v ImVec2, mn ImVec2, mx ImVec2)

@[c: 'igImLerp_Vec2Float']
fn im_lerp_vec2_float(p_out &ImVec2, a ImVec2, b ImVec2, t f32)

@[c: 'igImLerp_Vec2Vec2']
fn im_lerp_vec2_vec2(p_out &ImVec2, a ImVec2, b ImVec2, t ImVec2)

@[c: 'igImLerp_Vec4']
fn im_lerp_vec4(p_out &C.ImVec4, a C.ImVec4, b C.ImVec4, t f32)

@[c: 'igImSaturate']
fn im_saturate(f f32) f32

@[c: 'igImLengthSqr_Vec2']
fn im_length_sqr_vec2(lhs ImVec2) f32

@[c: 'igImLengthSqr_Vec4']
fn im_length_sqr_vec4(lhs C.ImVec4) f32

@[c: 'igImInvLength']
fn im_inv_length(lhs ImVec2, fail_value f32) f32

@[c: 'igImTrunc_Float']
fn im_trunc_float(f f32) f32

@[c: 'igImTrunc_Vec2']
fn im_trunc_vec2(p_out &ImVec2, v ImVec2)

@[c: 'igImFloor_Float']
fn im_floor_float(f f32) f32

@[c: 'igImFloor_Vec2']
fn im_floor_vec2(p_out &ImVec2, v ImVec2)

@[c: 'igImModPositive']
fn im_mod_positive(a int, b int) int

@[c: 'igImDot']
fn im_dot(a ImVec2, b ImVec2) f32

@[c: 'igImRotate']
fn im_rotate(p_out &ImVec2, v ImVec2, cos_a f32, sin_a f32)

@[c: 'igImLinearSweep']
fn im_linear_sweep(current f32, target f32, speed f32) f32

@[c: 'igImLinearRemapClamp']
fn im_linear_remap_clamp(s0 f32, s1 f32, d0 f32, d1 f32, x f32) f32

@[c: 'igImMul']
fn im_mul(p_out &ImVec2, lhs ImVec2, rhs ImVec2)

@[c: 'igImIsFloatAboveGuaranteedIntegerPrecision']
fn im_is_float_above_guaranteed_integer_precision(f f32) bool

@[c: 'igImExponentialMovingAverage']
fn im_exponential_moving_average(avg f32, sample f32, n int) f32

@[c: 'igImBezierCubicCalc']
fn im_bezier_cubic_calc(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, t f32)

@[c: 'igImBezierCubicClosestPoint']
fn im_bezier_cubic_closest_point(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, p ImVec2, num_segments int)

@[c: 'igImBezierCubicClosestPointCasteljau']
fn im_bezier_cubic_closest_point_casteljau(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, p ImVec2, tess_tol f32)

@[c: 'igImBezierQuadraticCalc']
fn im_bezier_quadratic_calc(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, t f32)

@[c: 'igImLineClosestPoint']
fn im_line_closest_point(p_out &ImVec2, a ImVec2, b ImVec2, p ImVec2)

@[c: 'igImTriangleContainsPoint']
fn im_triangle_contains_point(a ImVec2, b ImVec2, c ImVec2, p ImVec2) bool

@[c: 'igImTriangleClosestPoint']
fn im_triangle_closest_point(p_out &ImVec2, a ImVec2, b ImVec2, c ImVec2, p ImVec2)

@[c: 'igImTriangleBarycentricCoords']
fn im_triangle_barycentric_coords(a ImVec2, b ImVec2, c ImVec2, p ImVec2, out_u &f32, out_v &f32, out_w &f32)

@[c: 'igImTriangleArea']
fn im_triangle_area(a ImVec2, b ImVec2, c ImVec2) f32

@[c: 'igImTriangleIsClockwise']
fn im_triangle_is_clockwise(a ImVec2, b ImVec2, c ImVec2) bool

@[c: 'ImVec1_ImVec1_Nil']
fn im_vec1_im_vec1_nil() &ImVec1

@[c: 'ImVec1_ImVec1_Nil_Construct']
fn im_vec1_im_vec1_nil_construct(self &ImVec1)

@[c: 'ImVec1_destroy']
fn im_vec1_destroy(self &ImVec1)

@[c: 'ImVec1_ImVec1_Float']
fn im_vec1_im_vec1_float(_x f32) &ImVec1

@[c: 'ImVec1_ImVec1_Float_Construct']
fn im_vec1_im_vec1_float_construct(self &ImVec1, _x f32)

@[c: 'ImVec2ih_ImVec2ih_Nil']
fn im_vec2ih_im_vec2ih_nil() &ImVec2ih

@[c: 'ImVec2ih_ImVec2ih_Nil_Construct']
fn im_vec2ih_im_vec2ih_nil_construct(self &ImVec2ih)

@[c: 'ImVec2ih_destroy']
fn im_vec2ih_destroy(self &ImVec2ih)

@[c: 'ImVec2ih_ImVec2ih_short']
fn im_vec2ih_im_vec2ih_short(_x i16, _y i16) &ImVec2ih

@[c: 'ImVec2ih_ImVec2ih_short_Construct']
fn im_vec2ih_im_vec2ih_short_construct(self &ImVec2ih, _x i16, _y i16)

@[c: 'ImVec2ih_ImVec2ih_Vec2']
fn im_vec2ih_im_vec2ih_vec2(rhs ImVec2) &ImVec2ih

@[c: 'ImVec2ih_ImVec2ih_Vec2_Construct']
fn im_vec2ih_im_vec2ih_vec2_construct(self &ImVec2ih, rhs ImVec2)

@[c: 'ImRect_ImRect_Nil']
fn im_rect_im_rect_nil() &C.ImRect

@[c: 'ImRect_ImRect_Nil_Construct']
fn im_rect_im_rect_nil_construct(self &C.ImRect)

@[c: 'ImRect_destroy']
fn im_rect_destroy(self &C.ImRect)

@[c: 'ImRect_ImRect_Vec2']
fn im_rect_im_rect_vec2(min ImVec2, max ImVec2) &C.ImRect

@[c: 'ImRect_ImRect_Vec2_Construct']
fn im_rect_im_rect_vec2_construct(self &C.ImRect, min ImVec2, max ImVec2)

@[c: 'ImRect_ImRect_Vec4']
fn im_rect_im_rect_vec4(v C.ImVec4) &C.ImRect

@[c: 'ImRect_ImRect_Vec4_Construct']
fn im_rect_im_rect_vec4_construct(self &C.ImRect, v C.ImVec4)

@[c: 'ImRect_ImRect_Float']
fn im_rect_im_rect_float(x1 f32, y1 f32, x2 f32, y2 f32) &C.ImRect

@[c: 'ImRect_ImRect_Float_Construct']
fn im_rect_im_rect_float_construct(self &C.ImRect, x1 f32, y1 f32, x2 f32, y2 f32)

@[c: 'ImRect_GetCenter']
fn im_rect_get_center(p_out &ImVec2, self &C.ImRect)

@[c: 'ImRect_GetSize']
fn im_rect_get_size(p_out &ImVec2, self &C.ImRect)

@[c: 'ImRect_GetWidth']
fn im_rect_get_width(self &C.ImRect) f32

@[c: 'ImRect_GetHeight']
fn im_rect_get_height(self &C.ImRect) f32

@[c: 'ImRect_GetArea']
fn im_rect_get_area(self &C.ImRect) f32

@[c: 'ImRect_GetTL']
fn im_rect_get_tl(p_out &ImVec2, self &C.ImRect)

@[c: 'ImRect_GetTR']
fn im_rect_get_tr(p_out &ImVec2, self &C.ImRect)

@[c: 'ImRect_GetBL']
fn im_rect_get_bl(p_out &ImVec2, self &C.ImRect)

@[c: 'ImRect_GetBR']
fn im_rect_get_br(p_out &ImVec2, self &C.ImRect)

@[c: 'ImRect_Contains_Vec2']
fn im_rect_contains_vec2(self &C.ImRect, p ImVec2) bool

@[c: 'ImRect_Contains_Rect']
fn im_rect_contains_rect(self &C.ImRect, r C.ImRect) bool

@[c: 'ImRect_ContainsWithPad']
fn im_rect_contains_with_pad(self &C.ImRect, p ImVec2, pad ImVec2) bool

@[c: 'ImRect_Overlaps']
fn im_rect_overlaps(self &C.ImRect, r C.ImRect) bool

@[c: 'ImRect_Add_Vec2']
fn im_rect_add_vec2(self &C.ImRect, p ImVec2)

@[c: 'ImRect_Add_Rect']
fn im_rect_add_rect(self &C.ImRect, r C.ImRect)

@[c: 'ImRect_Expand_Float']
fn im_rect_expand_float(self &C.ImRect, amount f32)

@[c: 'ImRect_Expand_Vec2']
fn im_rect_expand_vec2(self &C.ImRect, amount ImVec2)

@[c: 'ImRect_Translate']
fn im_rect_translate(self &C.ImRect, d ImVec2)

@[c: 'ImRect_TranslateX']
fn im_rect_translate_x(self &C.ImRect, dx f32)

@[c: 'ImRect_TranslateY']
fn im_rect_translate_y(self &C.ImRect, dy f32)

@[c: 'ImRect_ClipWith']
fn im_rect_clip_with(self &C.ImRect, r C.ImRect)

@[c: 'ImRect_ClipWithFull']
fn im_rect_clip_with_full(self &C.ImRect, r C.ImRect)

@[c: 'ImRect_Floor']
fn im_rect_floor(self &C.ImRect)

@[c: 'ImRect_IsInverted']
fn im_rect_is_inverted(self &C.ImRect) bool

@[c: 'ImRect_ToVec4']
fn im_rect_to_vec4(p_out &C.ImVec4, self &C.ImRect)

@[c: 'igImBitArrayGetStorageSizeInBytes']
fn im_bit_array_get_storage_size_in_bytes(bitcount int) usize

@[c: 'igImBitArrayClearAllBits']
fn im_bit_array_clear_all_bits(arr &ImU32, bitcount int)

@[c: 'igImBitArrayTestBit']
fn im_bit_array_test_bit(arr &ImU32, n int) bool

@[c: 'igImBitArrayClearBit']
fn im_bit_array_clear_bit(arr &ImU32, n int)

@[c: 'igImBitArraySetBit']
fn im_bit_array_set_bit(arr &ImU32, n int)

@[c: 'igImBitArraySetBitRange']
fn im_bit_array_set_bit_range(arr &ImU32, n int, n2 int)

@[c: 'ImBitVector_Create']
fn im_bit_vector_create(self &C.ImBitVector, sz int)

@[c: 'ImBitVector_Clear']
fn im_bit_vector_clear(self &C.ImBitVector)

@[c: 'ImBitVector_TestBit']
fn im_bit_vector_test_bit(self &C.ImBitVector, n int) bool

@[c: 'ImBitVector_SetBit']
fn im_bit_vector_set_bit(self &C.ImBitVector, n int)

@[c: 'ImBitVector_ClearBit']
fn im_bit_vector_clear_bit(self &C.ImBitVector, n int)

@[c: 'ImGuiTextIndex_clear']
fn text_index_clear(self &TextIndex)

@[c: 'ImGuiTextIndex_size']
fn text_index_size(self &TextIndex) int

@[c: 'ImGuiTextIndex_get_line_begin']
fn text_index_get_line_begin(self &TextIndex, base &i8, n int) &i8

@[c: 'ImGuiTextIndex_get_line_end']
fn text_index_get_line_end(self &TextIndex, base &i8, n int) &i8

@[c: 'ImGuiTextIndex_append']
fn text_index_append(self &TextIndex, base &i8, old_size int, new_size int)

@[c: 'igImLowerBound']
fn im_lower_bound(in_begin &StoragePair, in_end &StoragePair, key ID) &StoragePair

@[c: 'ImDrawListSharedData_ImDrawListSharedData']
fn im_draw_list_shared_data_im_draw_list_shared_data() &ImDrawListSharedData

@[c: 'ImDrawListSharedData_ImDrawListSharedData_Construct']
fn im_draw_list_shared_data_im_draw_list_shared_data_construct(self &ImDrawListSharedData)

@[c: 'ImDrawListSharedData_destroy']
fn im_draw_list_shared_data_destroy(self &ImDrawListSharedData)

@[c: 'ImDrawListSharedData_SetCircleTessellationMaxError']
fn im_draw_list_shared_data_set_circle_tessellation_max_error(self &ImDrawListSharedData, max_error f32)

@[c: 'ImDrawDataBuilder_ImDrawDataBuilder']
fn im_draw_data_builder_im_draw_data_builder() &ImDrawDataBuilder

@[c: 'ImDrawDataBuilder_ImDrawDataBuilder_Construct']
fn im_draw_data_builder_im_draw_data_builder_construct(self &ImDrawDataBuilder)

@[c: 'ImDrawDataBuilder_destroy']
fn im_draw_data_builder_destroy(self &ImDrawDataBuilder)

@[c: 'ImGuiStyleVarInfo_GetVarPtr']
fn style_var_info_get_var_ptr(self &StyleVarInfo, parent voidptr) voidptr

@[c: 'ImGuiStyleMod_ImGuiStyleMod_Int']
fn style_mod_im_gui_style_mod_int(idx StyleVar, v int) &StyleMod

@[c: 'ImGuiStyleMod_ImGuiStyleMod_Int_Construct']
fn style_mod_im_gui_style_mod_int_construct(self &StyleMod, idx StyleVar, v int)

@[c: 'ImGuiStyleMod_destroy']
fn style_mod_destroy(self &StyleMod)

@[c: 'ImGuiStyleMod_ImGuiStyleMod_Float']
fn style_mod_im_gui_style_mod_float(idx StyleVar, v f32) &StyleMod

@[c: 'ImGuiStyleMod_ImGuiStyleMod_Float_Construct']
fn style_mod_im_gui_style_mod_float_construct(self &StyleMod, idx StyleVar, v f32)

@[c: 'ImGuiStyleMod_ImGuiStyleMod_Vec2']
fn style_mod_im_gui_style_mod_vec2(idx StyleVar, v ImVec2) &StyleMod

@[c: 'ImGuiStyleMod_ImGuiStyleMod_Vec2_Construct']
fn style_mod_im_gui_style_mod_vec2_construct(self &StyleMod, idx StyleVar, v ImVec2)

@[c: 'ImGuiComboPreviewData_ImGuiComboPreviewData']
fn combo_preview_data_im_gui_combo_preview_data() &ComboPreviewData

@[c: 'ImGuiComboPreviewData_ImGuiComboPreviewData_Construct']
fn combo_preview_data_im_gui_combo_preview_data_construct(self &ComboPreviewData)

@[c: 'ImGuiComboPreviewData_destroy']
fn combo_preview_data_destroy(self &ComboPreviewData)

@[c: 'ImGuiMenuColumns_ImGuiMenuColumns']
fn menu_columns_im_gui_menu_columns() &MenuColumns

@[c: 'ImGuiMenuColumns_ImGuiMenuColumns_Construct']
fn menu_columns_im_gui_menu_columns_construct(self &MenuColumns)

@[c: 'ImGuiMenuColumns_destroy']
fn menu_columns_destroy(self &MenuColumns)

@[c: 'ImGuiMenuColumns_Update']
fn menu_columns_update(self &MenuColumns, spacing f32, window_reappearing bool)

@[c: 'ImGuiMenuColumns_DeclColumns']
fn menu_columns_decl_columns(self &MenuColumns, w_icon f32, w_label f32, w_shortcut f32, w_mark f32) f32

@[c: 'ImGuiMenuColumns_CalcNextTotalWidth']
fn menu_columns_calc_next_total_width(self &MenuColumns, update_offsets bool)

@[c: 'ImGuiInputTextDeactivatedState_ImGuiInputTextDeactivatedState']
fn input_text_deactivated_state_im_gui_input_text_deactivated_state() &InputTextDeactivatedState

@[c: 'ImGuiInputTextDeactivatedState_ImGuiInputTextDeactivatedState_Construct']
fn input_text_deactivated_state_im_gui_input_text_deactivated_state_construct(self &InputTextDeactivatedState)

@[c: 'ImGuiInputTextDeactivatedState_destroy']
fn input_text_deactivated_state_destroy(self &InputTextDeactivatedState)

@[c: 'ImGuiInputTextDeactivatedState_ClearFreeMemory']
fn input_text_deactivated_state_clear_free_memory(self &InputTextDeactivatedState)

@[c: 'ImGuiInputTextState_ImGuiInputTextState']
fn input_text_state_im_gui_input_text_state() &InputTextState

@[c: 'ImGuiInputTextState_ImGuiInputTextState_Construct']
fn input_text_state_im_gui_input_text_state_construct(self &InputTextState)

@[c: 'ImGuiInputTextState_destroy']
fn input_text_state_destroy(self &InputTextState)

@[c: 'ImGuiInputTextState_ClearText']
fn input_text_state_clear_text(self &InputTextState)

@[c: 'ImGuiInputTextState_ClearFreeMemory']
fn input_text_state_clear_free_memory(self &InputTextState)

@[c: 'ImGuiInputTextState_OnKeyPressed']
fn input_text_state_on_key_pressed(self &InputTextState, key int)

@[c: 'ImGuiInputTextState_OnCharPressed']
fn input_text_state_on_char_pressed(self &InputTextState, c u32)

@[c: 'ImGuiInputTextState_CursorAnimReset']
fn input_text_state_cursor_anim_reset(self &InputTextState)

@[c: 'ImGuiInputTextState_CursorClamp']
fn input_text_state_cursor_clamp(self &InputTextState)

@[c: 'ImGuiInputTextState_HasSelection']
fn input_text_state_has_selection(self &InputTextState) bool

@[c: 'ImGuiInputTextState_ClearSelection']
fn input_text_state_clear_selection(self &InputTextState)

@[c: 'ImGuiInputTextState_GetCursorPos']
fn input_text_state_get_cursor_pos(self &InputTextState) int

@[c: 'ImGuiInputTextState_GetSelectionStart']
fn input_text_state_get_selection_start(self &InputTextState) int

@[c: 'ImGuiInputTextState_GetSelectionEnd']
fn input_text_state_get_selection_end(self &InputTextState) int

@[c: 'ImGuiInputTextState_SelectAll']
fn input_text_state_select_all(self &InputTextState)

@[c: 'ImGuiInputTextState_ReloadUserBufAndSelectAll']
fn input_text_state_reload_user_buf_and_select_all(self &InputTextState)

@[c: 'ImGuiInputTextState_ReloadUserBufAndKeepSelection']
fn input_text_state_reload_user_buf_and_keep_selection(self &InputTextState)

@[c: 'ImGuiInputTextState_ReloadUserBufAndMoveToEnd']
fn input_text_state_reload_user_buf_and_move_to_end(self &InputTextState)

@[c: 'ImGuiNextWindowData_ImGuiNextWindowData']
fn next_window_data_im_gui_next_window_data() &NextWindowData

@[c: 'ImGuiNextWindowData_ImGuiNextWindowData_Construct']
fn next_window_data_im_gui_next_window_data_construct(self &NextWindowData)

@[c: 'ImGuiNextWindowData_destroy']
fn next_window_data_destroy(self &NextWindowData)

@[c: 'ImGuiNextWindowData_ClearFlags']
fn next_window_data_clear_flags(self &NextWindowData)

@[c: 'ImGuiNextItemData_ImGuiNextItemData']
fn next_item_data_im_gui_next_item_data() &NextItemData

@[c: 'ImGuiNextItemData_ImGuiNextItemData_Construct']
fn next_item_data_im_gui_next_item_data_construct(self &NextItemData)

@[c: 'ImGuiNextItemData_destroy']
fn next_item_data_destroy(self &NextItemData)

@[c: 'ImGuiNextItemData_ClearFlags']
fn next_item_data_clear_flags(self &NextItemData)

@[c: 'ImGuiLastItemData_ImGuiLastItemData']
fn last_item_data_im_gui_last_item_data() &LastItemData

@[c: 'ImGuiLastItemData_ImGuiLastItemData_Construct']
fn last_item_data_im_gui_last_item_data_construct(self &LastItemData)

@[c: 'ImGuiLastItemData_destroy']
fn last_item_data_destroy(self &LastItemData)

@[c: 'ImGuiErrorRecoveryState_ImGuiErrorRecoveryState']
fn error_recovery_state_im_gui_error_recovery_state() &ErrorRecoveryState

@[c: 'ImGuiErrorRecoveryState_ImGuiErrorRecoveryState_Construct']
fn error_recovery_state_im_gui_error_recovery_state_construct(self &ErrorRecoveryState)

@[c: 'ImGuiErrorRecoveryState_destroy']
fn error_recovery_state_destroy(self &ErrorRecoveryState)

@[c: 'ImGuiPtrOrIndex_ImGuiPtrOrIndex_Ptr']
fn ptr_or_index_im_gui_ptr_or_index_ptr(ptr voidptr) &PtrOrIndex

@[c: 'ImGuiPtrOrIndex_ImGuiPtrOrIndex_Ptr_Construct']
fn ptr_or_index_im_gui_ptr_or_index_ptr_construct(self &PtrOrIndex, ptr voidptr)

@[c: 'ImGuiPtrOrIndex_destroy']
fn ptr_or_index_destroy(self &PtrOrIndex)

@[c: 'ImGuiPtrOrIndex_ImGuiPtrOrIndex_Int']
fn ptr_or_index_im_gui_ptr_or_index_int(index int) &PtrOrIndex

@[c: 'ImGuiPtrOrIndex_ImGuiPtrOrIndex_Int_Construct']
fn ptr_or_index_im_gui_ptr_or_index_int_construct(self &PtrOrIndex, index int)

@[c: 'ImGuiPopupData_ImGuiPopupData']
fn popup_data_im_gui_popup_data() &PopupData

@[c: 'ImGuiPopupData_ImGuiPopupData_Construct']
fn popup_data_im_gui_popup_data_construct(self &PopupData)

@[c: 'ImGuiPopupData_destroy']
fn popup_data_destroy(self &PopupData)

@[c: 'ImGuiInputEvent_ImGuiInputEvent']
fn input_event_im_gui_input_event() &C.ImGuiInputEvent

@[c: 'ImGuiInputEvent_ImGuiInputEvent_Construct']
fn input_event_im_gui_input_event_construct(self &C.ImGuiInputEvent)

@[c: 'ImGuiInputEvent_destroy']
fn input_event_destroy(self &C.ImGuiInputEvent)

@[c: 'ImGuiKeyRoutingData_ImGuiKeyRoutingData']
fn key_routing_data_im_gui_key_routing_data() &KeyRoutingData

@[c: 'ImGuiKeyRoutingData_ImGuiKeyRoutingData_Construct']
fn key_routing_data_im_gui_key_routing_data_construct(self &KeyRoutingData)

@[c: 'ImGuiKeyRoutingData_destroy']
fn key_routing_data_destroy(self &KeyRoutingData)

@[c: 'ImGuiKeyRoutingTable_ImGuiKeyRoutingTable']
fn key_routing_table_im_gui_key_routing_table() &KeyRoutingTable

@[c: 'ImGuiKeyRoutingTable_ImGuiKeyRoutingTable_Construct']
fn key_routing_table_im_gui_key_routing_table_construct(self &KeyRoutingTable)

@[c: 'ImGuiKeyRoutingTable_destroy']
fn key_routing_table_destroy(self &KeyRoutingTable)

@[c: 'ImGuiKeyRoutingTable_Clear']
fn key_routing_table_clear(self &KeyRoutingTable)

@[c: 'ImGuiKeyOwnerData_ImGuiKeyOwnerData']
fn key_owner_data_im_gui_key_owner_data() &KeyOwnerData

@[c: 'ImGuiKeyOwnerData_ImGuiKeyOwnerData_Construct']
fn key_owner_data_im_gui_key_owner_data_construct(self &KeyOwnerData)

@[c: 'ImGuiKeyOwnerData_destroy']
fn key_owner_data_destroy(self &KeyOwnerData)

@[c: 'ImGuiListClipperRange_FromIndices']
fn list_clipper_range_from_indices(min int, max int) ListClipperRange

@[c: 'ImGuiListClipperRange_FromPositions']
fn list_clipper_range_from_positions(y1 f32, y2 f32, off_min int, off_max int) ListClipperRange

@[c: 'ImGuiListClipperData_ImGuiListClipperData']
fn list_clipper_data_im_gui_list_clipper_data() &ListClipperData

@[c: 'ImGuiListClipperData_ImGuiListClipperData_Construct']
fn list_clipper_data_im_gui_list_clipper_data_construct(self &ListClipperData)

@[c: 'ImGuiListClipperData_destroy']
fn list_clipper_data_destroy(self &ListClipperData)

@[c: 'ImGuiListClipperData_Reset']
fn list_clipper_data_reset(self &ListClipperData, clipper &ListClipper)

@[c: 'ImGuiNavItemData_ImGuiNavItemData']
fn nav_item_data_im_gui_nav_item_data() &NavItemData

@[c: 'ImGuiNavItemData_ImGuiNavItemData_Construct']
fn nav_item_data_im_gui_nav_item_data_construct(self &NavItemData)

@[c: 'ImGuiNavItemData_destroy']
fn nav_item_data_destroy(self &NavItemData)

@[c: 'ImGuiNavItemData_Clear']
fn nav_item_data_clear(self &NavItemData)

@[c: 'ImGuiTypingSelectState_ImGuiTypingSelectState']
fn typing_select_state_im_gui_typing_select_state() &TypingSelectState

@[c: 'ImGuiTypingSelectState_ImGuiTypingSelectState_Construct']
fn typing_select_state_im_gui_typing_select_state_construct(self &TypingSelectState)

@[c: 'ImGuiTypingSelectState_destroy']
fn typing_select_state_destroy(self &TypingSelectState)

@[c: 'ImGuiTypingSelectState_Clear']
fn typing_select_state_clear(self &TypingSelectState)

@[c: 'ImGuiOldColumnData_ImGuiOldColumnData']
fn old_column_data_im_gui_old_column_data() &OldColumnData

@[c: 'ImGuiOldColumnData_ImGuiOldColumnData_Construct']
fn old_column_data_im_gui_old_column_data_construct(self &OldColumnData)

@[c: 'ImGuiOldColumnData_destroy']
fn old_column_data_destroy(self &OldColumnData)

@[c: 'ImGuiOldColumns_ImGuiOldColumns']
fn old_columns_im_gui_old_columns() &OldColumns

@[c: 'ImGuiOldColumns_ImGuiOldColumns_Construct']
fn old_columns_im_gui_old_columns_construct(self &OldColumns)

@[c: 'ImGuiOldColumns_destroy']
fn old_columns_destroy(self &OldColumns)

@[c: 'ImGuiBoxSelectState_ImGuiBoxSelectState']
fn box_select_state_im_gui_box_select_state() &BoxSelectState

@[c: 'ImGuiBoxSelectState_ImGuiBoxSelectState_Construct']
fn box_select_state_im_gui_box_select_state_construct(self &BoxSelectState)

@[c: 'ImGuiBoxSelectState_destroy']
fn box_select_state_destroy(self &BoxSelectState)

@[c: 'ImGuiMultiSelectTempData_ImGuiMultiSelectTempData']
fn multi_select_temp_data_im_gui_multi_select_temp_data() &MultiSelectTempData

@[c: 'ImGuiMultiSelectTempData_ImGuiMultiSelectTempData_Construct']
fn multi_select_temp_data_im_gui_multi_select_temp_data_construct(self &MultiSelectTempData)

@[c: 'ImGuiMultiSelectTempData_destroy']
fn multi_select_temp_data_destroy(self &MultiSelectTempData)

@[c: 'ImGuiMultiSelectTempData_Clear']
fn multi_select_temp_data_clear(self &MultiSelectTempData)

@[c: 'ImGuiMultiSelectTempData_ClearIO']
fn multi_select_temp_data_clear_io(self &MultiSelectTempData)

@[c: 'ImGuiMultiSelectState_ImGuiMultiSelectState']
fn multi_select_state_im_gui_multi_select_state() &MultiSelectState

@[c: 'ImGuiMultiSelectState_ImGuiMultiSelectState_Construct']
fn multi_select_state_im_gui_multi_select_state_construct(self &MultiSelectState)

@[c: 'ImGuiMultiSelectState_destroy']
fn multi_select_state_destroy(self &MultiSelectState)

@[c: 'ImGuiDockNode_ImGuiDockNode']
fn dock_node_im_gui_dock_node(id ID) &DockNode

@[c: 'ImGuiDockNode_ImGuiDockNode_Construct']
fn dock_node_im_gui_dock_node_construct(self &DockNode, id ID)

@[c: 'ImGuiDockNode_destroy']
fn dock_node_destroy(self &DockNode)

@[c: 'ImGuiDockNode_IsRootNode']
fn dock_node_is_root_node(self &DockNode) bool

@[c: 'ImGuiDockNode_IsDockSpace']
fn dock_node_is_dock_space(self &DockNode) bool

@[c: 'ImGuiDockNode_IsFloatingNode']
fn dock_node_is_floating_node(self &DockNode) bool

@[c: 'ImGuiDockNode_IsCentralNode']
fn dock_node_is_central_node(self &DockNode) bool

@[c: 'ImGuiDockNode_IsHiddenTabBar']
fn dock_node_is_hidden_tab_bar(self &DockNode) bool

@[c: 'ImGuiDockNode_IsNoTabBar']
fn dock_node_is_no_tab_bar(self &DockNode) bool

@[c: 'ImGuiDockNode_IsSplitNode']
fn dock_node_is_split_node(self &DockNode) bool

@[c: 'ImGuiDockNode_IsLeafNode']
fn dock_node_is_leaf_node(self &DockNode) bool

@[c: 'ImGuiDockNode_IsEmpty']
fn dock_node_is_empty(self &DockNode) bool

@[c: 'ImGuiDockNode_Rect']
fn dock_node_rect(p_out &C.ImRect, self &DockNode)

@[c: 'ImGuiDockNode_SetLocalFlags']
fn dock_node_set_local_flags(self &DockNode, flags DockNodeFlags)

@[c: 'ImGuiDockNode_UpdateMergedFlags']
fn dock_node_update_merged_flags(self &DockNode)

@[c: 'ImGuiDockContext_ImGuiDockContext']
fn dock_context_im_gui_dock_context() &DockContext

@[c: 'ImGuiDockContext_ImGuiDockContext_Construct']
fn dock_context_im_gui_dock_context_construct(self &DockContext)

@[c: 'ImGuiDockContext_destroy']
fn dock_context_destroy(self &DockContext)

@[c: 'ImGuiViewportP_ImGuiViewportP']
fn viewport_p_im_gui_viewport_p() &ViewportP

@[c: 'ImGuiViewportP_ImGuiViewportP_Construct']
fn viewport_p_im_gui_viewport_p_construct(self &ViewportP)

@[c: 'ImGuiViewportP_destroy']
fn viewport_p_destroy(self &ViewportP)

@[c: 'ImGuiViewportP_ClearRequestFlags']
fn viewport_p_clear_request_flags(self &ViewportP)

@[c: 'ImGuiViewportP_CalcWorkRectPos']
fn viewport_p_calc_work_rect_pos(p_out &ImVec2, self &ViewportP, inset_min ImVec2)

@[c: 'ImGuiViewportP_CalcWorkRectSize']
fn viewport_p_calc_work_rect_size(p_out &ImVec2, self &ViewportP, inset_min ImVec2, inset_max ImVec2)

@[c: 'ImGuiViewportP_UpdateWorkRect']
fn viewport_p_update_work_rect(self &ViewportP)

@[c: 'ImGuiViewportP_GetMainRect']
fn viewport_p_get_main_rect(p_out &C.ImRect, self &ViewportP)

@[c: 'ImGuiViewportP_GetWorkRect']
fn viewport_p_get_work_rect(p_out &C.ImRect, self &ViewportP)

@[c: 'ImGuiViewportP_GetBuildWorkRect']
fn viewport_p_get_build_work_rect(p_out &C.ImRect, self &ViewportP)

@[c: 'ImGuiWindowSettings_ImGuiWindowSettings']
fn window_settings_im_gui_window_settings() &WindowSettings

@[c: 'ImGuiWindowSettings_ImGuiWindowSettings_Construct']
fn window_settings_im_gui_window_settings_construct(self &WindowSettings)

@[c: 'ImGuiWindowSettings_destroy']
fn window_settings_destroy(self &WindowSettings)

@[c: 'ImGuiWindowSettings_GetName']
fn window_settings_get_name(self &WindowSettings) &i8

@[c: 'ImGuiSettingsHandler_ImGuiSettingsHandler']
fn settings_handler_im_gui_settings_handler() &SettingsHandler

@[c: 'ImGuiSettingsHandler_ImGuiSettingsHandler_Construct']
fn settings_handler_im_gui_settings_handler_construct(self &SettingsHandler)

@[c: 'ImGuiSettingsHandler_destroy']
fn settings_handler_destroy(self &SettingsHandler)

@[c: 'ImGuiDebugAllocInfo_ImGuiDebugAllocInfo']
fn debug_alloc_info_im_gui_debug_alloc_info() &DebugAllocInfo

@[c: 'ImGuiDebugAllocInfo_ImGuiDebugAllocInfo_Construct']
fn debug_alloc_info_im_gui_debug_alloc_info_construct(self &DebugAllocInfo)

@[c: 'ImGuiDebugAllocInfo_destroy']
fn debug_alloc_info_destroy(self &DebugAllocInfo)

@[c: 'ImGuiStackLevelInfo_ImGuiStackLevelInfo']
fn stack_level_info_im_gui_stack_level_info() &StackLevelInfo

@[c: 'ImGuiStackLevelInfo_ImGuiStackLevelInfo_Construct']
fn stack_level_info_im_gui_stack_level_info_construct(self &StackLevelInfo)

@[c: 'ImGuiStackLevelInfo_destroy']
fn stack_level_info_destroy(self &StackLevelInfo)

@[c: 'ImGuiIDStackTool_ImGuiIDStackTool']
fn ids_tack_tool_im_gui_ids_tack_tool() &C.ImGuiIDStackTool

@[c: 'ImGuiIDStackTool_ImGuiIDStackTool_Construct']
fn ids_tack_tool_im_gui_ids_tack_tool_construct(self &C.ImGuiIDStackTool)

@[c: 'ImGuiIDStackTool_destroy']
fn ids_tack_tool_destroy(self &C.ImGuiIDStackTool)

@[c: 'ImGuiContextHook_ImGuiContextHook']
fn context_hook_im_gui_context_hook() &ContextHook

@[c: 'ImGuiContextHook_ImGuiContextHook_Construct']
fn context_hook_im_gui_context_hook_construct(self &ContextHook)

@[c: 'ImGuiContextHook_destroy']
fn context_hook_destroy(self &ContextHook)

@[c: 'ImGuiContext_ImGuiContext']
fn context_im_gui_context(shared_font_atlas &ImFontAtlas) &Context

@[c: 'ImGuiContext_ImGuiContext_Construct']
fn context_im_gui_context_construct(self &Context, shared_font_atlas &ImFontAtlas)

@[c: 'ImGuiContext_destroy']
fn context_destroy(self &Context)

@[c: 'ImGuiWindow_ImGuiWindow']
fn window_im_gui_window(context &Context, name &i8) &Window

@[c: 'ImGuiWindow_ImGuiWindow_Construct']
fn window_im_gui_window_construct(self &Window, context &Context, name &i8)

@[c: 'ImGuiWindow_destroy']
fn window_destroy(self &Window)

@[c: 'ImGuiWindow_GetID_Str']
fn window_get_id_str(self &Window, str &i8, str_end &i8) ID

@[c: 'ImGuiWindow_GetID_Ptr']
fn window_get_id_ptr(self &Window, ptr voidptr) ID

@[c: 'ImGuiWindow_GetID_Int']
fn window_get_id_int(self &Window, n int) ID

@[c: 'ImGuiWindow_GetIDFromPos']
fn window_get_idf_rom_pos(self &Window, p_abs ImVec2) ID

@[c: 'ImGuiWindow_GetIDFromRectangle']
fn window_get_idf_rom_rectangle(self &Window, r_abs C.ImRect) ID

@[c: 'ImGuiWindow_Rect']
fn window_rect(p_out &C.ImRect, self &Window)

@[c: 'ImGuiWindow_CalcFontSize']
fn window_calc_font_size(self &Window) f32

@[c: 'ImGuiWindow_TitleBarRect']
fn window_title_bar_rect(p_out &C.ImRect, self &Window)

@[c: 'ImGuiWindow_MenuBarRect']
fn window_menu_bar_rect(p_out &C.ImRect, self &Window)

@[c: 'ImGuiTabItem_ImGuiTabItem']
fn tab_item_im_gui_tab_item() &TabItem

@[c: 'ImGuiTabItem_ImGuiTabItem_Construct']
fn tab_item_im_gui_tab_item_construct(self &TabItem)

@[c: 'ImGuiTabItem_destroy']
fn tab_item_destroy(self &TabItem)

@[c: 'ImGuiTabBar_ImGuiTabBar']
fn tab_bar_im_gui_tab_bar() &C.ImGuiTabBar

@[c: 'ImGuiTabBar_ImGuiTabBar_Construct']
fn tab_bar_im_gui_tab_bar_construct(self &C.ImGuiTabBar)

@[c: 'ImGuiTabBar_destroy']
fn tab_bar_destroy(self &C.ImGuiTabBar)

@[c: 'ImGuiTableColumn_ImGuiTableColumn']
fn table_column_im_gui_table_column() &TableColumn

@[c: 'ImGuiTableColumn_ImGuiTableColumn_Construct']
fn table_column_im_gui_table_column_construct(self &TableColumn)

@[c: 'ImGuiTableColumn_destroy']
fn table_column_destroy(self &TableColumn)

@[c: 'ImGuiTableInstanceData_ImGuiTableInstanceData']
fn table_instance_data_im_gui_table_instance_data() &TableInstanceData

@[c: 'ImGuiTableInstanceData_ImGuiTableInstanceData_Construct']
fn table_instance_data_im_gui_table_instance_data_construct(self &TableInstanceData)

@[c: 'ImGuiTableInstanceData_destroy']
fn table_instance_data_destroy(self &TableInstanceData)

@[c: 'ImGuiTable_ImGuiTable']
fn table_im_gui_table() &Table

@[c: 'ImGuiTable_ImGuiTable_Construct']
fn table_im_gui_table_construct(self &Table)

@[c: 'ImGuiTable_destroy']
fn table_destroy(self &Table)

@[c: 'ImGuiTableTempData_ImGuiTableTempData']
fn table_temp_data_im_gui_table_temp_data() &TableTempData

@[c: 'ImGuiTableTempData_ImGuiTableTempData_Construct']
fn table_temp_data_im_gui_table_temp_data_construct(self &TableTempData)

@[c: 'ImGuiTableTempData_destroy']
fn table_temp_data_destroy(self &TableTempData)

@[c: 'ImGuiTableColumnSettings_ImGuiTableColumnSettings']
fn table_column_settings_im_gui_table_column_settings() &TableColumnSettings

@[c: 'ImGuiTableColumnSettings_ImGuiTableColumnSettings_Construct']
fn table_column_settings_im_gui_table_column_settings_construct(self &TableColumnSettings)

@[c: 'ImGuiTableColumnSettings_destroy']
fn table_column_settings_destroy(self &TableColumnSettings)

@[c: 'ImGuiTableSettings_ImGuiTableSettings']
fn table_settings_im_gui_table_settings() &TableSettings

@[c: 'ImGuiTableSettings_ImGuiTableSettings_Construct']
fn table_settings_im_gui_table_settings_construct(self &TableSettings)

@[c: 'ImGuiTableSettings_destroy']
fn table_settings_destroy(self &TableSettings)

@[c: 'ImGuiTableSettings_GetColumnSettings']
fn table_settings_get_column_settings(self &TableSettings) &TableColumnSettings

@[c: 'igGetIO_ContextPtr']
fn get_io_context_ptr(ctx &Context) &IO

@[c: 'igGetPlatformIO_ContextPtr']
fn get_platform_io_context_ptr(ctx &Context) &PlatformIO

@[c: 'igGetCurrentWindowRead']
fn get_current_window_read() &Window

@[c: 'igGetCurrentWindow']
fn get_current_window() &Window

@[c: 'igFindWindowByID']
fn find_window_by_id(id ID) &Window

@[c: 'igFindWindowByName']
fn find_window_by_name(name &i8) &Window

@[c: 'igUpdateWindowParentAndRootLinks']
fn update_window_parent_and_root_links(window &Window, flags WindowFlags, parent_window &Window)

@[c: 'igUpdateWindowSkipRefresh']
fn update_window_skip_refresh(window &Window)

@[c: 'igCalcWindowNextAutoFitSize']
fn calc_window_next_auto_fit_size(p_out &ImVec2, window &Window)

@[c: 'igIsWindowChildOf']
fn is_window_child_of(window &Window, potential_parent &Window, popup_hierarchy bool, dock_hierarchy bool) bool

@[c: 'igIsWindowWithinBeginStackOf']
fn is_window_within_begin_stack_of(window &Window, potential_parent &Window) bool

@[c: 'igIsWindowAbove']
fn is_window_above(potential_above &Window, potential_below &Window) bool

@[c: 'igIsWindowNavFocusable']
fn is_window_nav_focusable(window &Window) bool

@[c: 'igSetWindowPos_WindowPtr']
fn set_window_pos_window_ptr(window &Window, pos ImVec2, cond Cond)

@[c: 'igSetWindowSize_WindowPtr']
fn set_window_size_window_ptr(window &Window, size ImVec2, cond Cond)

@[c: 'igSetWindowCollapsed_WindowPtr']
fn set_window_collapsed_window_ptr(window &Window, collapsed bool, cond Cond)

@[c: 'igSetWindowHitTestHole']
fn set_window_hit_test_hole(window &Window, pos ImVec2, size ImVec2)

@[c: 'igSetWindowHiddenAndSkipItemsForCurrentFrame']
fn set_window_hidden_and_skip_items_for_current_frame(window &Window)

@[c: 'igSetWindowParentWindowForFocusRoute']
fn set_window_parent_window_for_focus_route(window &Window, parent_window &Window)

@[c: 'igWindowRectAbsToRel']
fn window_rect_abs_to_rel(p_out &C.ImRect, window &Window, r C.ImRect)

@[c: 'igWindowRectRelToAbs']
fn window_rect_rel_to_abs(p_out &C.ImRect, window &Window, r C.ImRect)

@[c: 'igWindowPosAbsToRel']
fn window_pos_abs_to_rel(p_out &ImVec2, window &Window, p ImVec2)

@[c: 'igWindowPosRelToAbs']
fn window_pos_rel_to_abs(p_out &ImVec2, window &Window, p ImVec2)

@[c: 'igFocusWindow']
fn focus_window(window &Window, flags FocusRequestFlags)

@[c: 'igFocusTopMostWindowUnderOne']
fn focus_top_most_window_under_one(under_this_window &Window, ignore_window &Window, filter_viewport &Viewport, flags FocusRequestFlags)

@[c: 'igBringWindowToFocusFront']
fn bring_window_to_focus_front(window &Window)

@[c: 'igBringWindowToDisplayFront']
fn bring_window_to_display_front(window &Window)

@[c: 'igBringWindowToDisplayBack']
fn bring_window_to_display_back(window &Window)

@[c: 'igBringWindowToDisplayBehind']
fn bring_window_to_display_behind(window &Window, above_window &Window)

@[c: 'igFindWindowDisplayIndex']
fn find_window_display_index(window &Window) int

@[c: 'igFindBottomMostVisibleWindowWithinBeginStack']
fn find_bottom_most_visible_window_within_begin_stack(window &Window) &Window

@[c: 'igSetNextWindowRefreshPolicy']
fn set_next_window_refresh_policy(flags WindowRefreshFlags)

@[c: 'igSetCurrentFont']
fn set_current_font(font &ImFont)

@[c: 'igGetDefaultFont']
fn get_default_font() &ImFont

@[c: 'igPushPasswordFont']
fn push_password_font()

@[c: 'igGetForegroundDrawList_WindowPtr']
fn get_foreground_draw_list_window_ptr(window &Window) &ImDrawList

@[c: 'igAddDrawListToDrawDataEx']
fn add_draw_list_to_draw_data_ex(draw_data &ImDrawData, out_list &ImVector_ImDrawListPtr, draw_list &ImDrawList)

@[c: 'igInitialize']
fn initialize()

@[c: 'igShutdown']
fn shutdown()

@[c: 'igUpdateInputEvents']
fn update_input_events(trickle_fast_inputs bool)

@[c: 'igUpdateHoveredWindowAndCaptureFlags']
fn update_hovered_window_and_capture_flags()

@[c: 'igFindHoveredWindowEx']
fn find_hovered_window_ex(pos ImVec2, find_first_and_in_any_viewport bool, out_hovered_window &&Window, out_hovered_window_under_moving_window &&Window)

@[c: 'igStartMouseMovingWindow']
fn start_mouse_moving_window(window &Window)

@[c: 'igStartMouseMovingWindowOrNode']
fn start_mouse_moving_window_or_node(window &Window, node &DockNode, undock bool)

@[c: 'igUpdateMouseMovingWindowNewFrame']
fn update_mouse_moving_window_new_frame()

@[c: 'igUpdateMouseMovingWindowEndFrame']
fn update_mouse_moving_window_end_frame()

@[c: 'igAddContextHook']
fn add_context_hook(context &Context, hook &ContextHook) ID

@[c: 'igRemoveContextHook']
fn remove_context_hook(context &Context, hook_to_remove ID)

@[c: 'igCallContextHooks']
fn call_context_hooks(context &Context, type_ ContextHookType)

@[c: 'igTranslateWindowsInViewport']
fn translate_windows_in_viewport(viewport &ViewportP, old_pos ImVec2, new_pos ImVec2, old_size ImVec2, new_size ImVec2)

@[c: 'igScaleWindowsInViewport']
fn scale_windows_in_viewport(viewport &ViewportP, scale f32)

@[c: 'igDestroyPlatformWindow']
fn destroy_platform_window(viewport &ViewportP)

@[c: 'igSetWindowViewport']
fn set_window_viewport(window &Window, viewport &ViewportP)

@[c: 'igSetCurrentViewport']
fn set_current_viewport(window &Window, viewport &ViewportP)

@[c: 'igGetViewportPlatformMonitor']
fn get_viewport_platform_monitor(viewport &Viewport) &PlatformMonitor

@[c: 'igFindHoveredViewportFromPlatformWindowStack']
fn find_hovered_viewport_from_platform_window_stack(mouse_platform_pos ImVec2) &ViewportP

@[c: 'igMarkIniSettingsDirty_Nil']
fn mark_ini_settings_dirty_nil()

@[c: 'igMarkIniSettingsDirty_WindowPtr']
fn mark_ini_settings_dirty_window_ptr(window &Window)

@[c: 'igClearIniSettings']
fn clear_ini_settings()

@[c: 'igAddSettingsHandler']
fn add_settings_handler(handler &SettingsHandler)

@[c: 'igRemoveSettingsHandler']
fn remove_settings_handler(type_name &i8)

@[c: 'igFindSettingsHandler']
fn find_settings_handler(type_name &i8) &SettingsHandler

@[c: 'igCreateNewWindowSettings']
fn create_new_window_settings(name &i8) &WindowSettings

@[c: 'igFindWindowSettingsByID']
fn find_window_settings_by_id(id ID) &WindowSettings

@[c: 'igFindWindowSettingsByWindow']
fn find_window_settings_by_window(window &Window) &WindowSettings

@[c: 'igClearWindowSettings']
fn clear_window_settings(name &i8)

@[c: 'igLocalizeRegisterEntries']
fn localize_register_entries(entries &C.ImGuiLocEntry, count int)

@[c: 'igLocalizeGetMsg']
fn localize_get_msg(key LocKey) &i8

@[c: 'igSetScrollX_WindowPtr']
fn set_scroll_x_window_ptr(window &Window, scroll_x f32)

@[c: 'igSetScrollY_WindowPtr']
fn set_scroll_y_window_ptr(window &Window, scroll_y f32)

@[c: 'igSetScrollFromPosX_WindowPtr']
fn set_scroll_from_pos_x_window_ptr(window &Window, local_x f32, center_x_ratio f32)

@[c: 'igSetScrollFromPosY_WindowPtr']
fn set_scroll_from_pos_y_window_ptr(window &Window, local_y f32, center_y_ratio f32)

@[c: 'igScrollToItem']
fn scroll_to_item(flags ScrollFlags)

@[c: 'igScrollToRect']
fn scroll_to_rect(window &Window, rect C.ImRect, flags ScrollFlags)

@[c: 'igScrollToRectEx']
fn scroll_to_rect_ex(p_out &ImVec2, window &Window, rect C.ImRect, flags ScrollFlags)

@[c: 'igScrollToBringRectIntoView']
fn scroll_to_bring_rect_into_view(window &Window, rect C.ImRect)

@[c: 'igGetItemStatusFlags']
fn get_item_status_flags() ItemStatusFlags

@[c: 'igGetItemFlags']
fn get_item_flags() ItemFlags

@[c: 'igGetActiveID']
fn get_active_id() ID

@[c: 'igGetFocusID']
fn get_focus_id() ID

@[c: 'igSetActiveID']
fn set_active_id(id ID, window &Window)

@[c: 'igSetFocusID']
fn set_focus_id(id ID, window &Window)

@[c: 'igClearActiveID']
fn clear_active_id()

@[c: 'igGetHoveredID']
fn get_hovered_id() ID

@[c: 'igSetHoveredID']
fn set_hovered_id(id ID)

@[c: 'igKeepAliveID']
fn keep_alive_id(id ID)

@[c: 'igMarkItemEdited']
fn mark_item_edited(id ID)

@[c: 'igPushOverrideID']
fn push_override_id(id ID)

@[c: 'igGetIDWithSeed_Str']
fn get_idw_ith_seed_str(str_id_begin &i8, str_id_end &i8, seed ID) ID

@[c: 'igGetIDWithSeed_Int']
fn get_idw_ith_seed_int(n int, seed ID) ID

@[c: 'igItemSize_Vec2']
fn item_size_vec2(size ImVec2, text_baseline_y f32)

@[c: 'igItemSize_Rect']
fn item_size_rect(bb C.ImRect, text_baseline_y f32)

@[c: 'igItemAdd']
fn item_add(bb C.ImRect, id ID, nav_bb &C.ImRect, extra_flags ItemFlags) bool

@[c: 'igItemHoverable']
fn item_hoverable(bb C.ImRect, id ID, item_flags ItemFlags) bool

@[c: 'igIsWindowContentHoverable']
fn is_window_content_hoverable(window &Window, flags HoveredFlags) bool

@[c: 'igIsClippedEx']
fn is_clipped_ex(bb C.ImRect, id ID) bool

@[c: 'igSetLastItemData']
fn set_last_item_data(item_id ID, item_flags ItemFlags, status_flags ItemStatusFlags, item_rect C.ImRect)

@[c: 'igCalcItemSize']
fn calc_item_size(p_out &ImVec2, size ImVec2, default_w f32, default_h f32)

@[c: 'igCalcWrapWidthForPos']
fn calc_wrap_width_for_pos(pos ImVec2, wrap_pos_x f32) f32

@[c: 'igPushMultiItemsWidths']
fn push_multi_items_widths(components int, width_full f32)

@[c: 'igShrinkWidths']
fn shrink_widths(items &ShrinkWidthItem, count int, width_excess f32)

@[c: 'igGetStyleVarInfo']
fn get_style_var_info(idx StyleVar) &StyleVarInfo

@[c: 'igBeginDisabledOverrideReenable']
fn begin_disabled_override_reenable()

@[c: 'igEndDisabledOverrideReenable']
fn end_disabled_override_reenable()

@[c: 'igLogBegin']
fn log_begin(flags LogFlags, auto_open_depth int)

@[c: 'igLogToBuffer']
fn log_to_buffer(auto_open_depth int)

@[c: 'igLogRenderedText']
fn log_rendered_text(ref_pos &ImVec2, text &i8, text_end &i8)

@[c: 'igLogSetNextTextDecoration']
fn log_set_next_text_decoration(prefix &i8, suffix &i8)

@[c: 'igBeginChildEx']
fn begin_child_ex(name &i8, id ID, size_arg ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c: 'igBeginPopupEx']
fn begin_popup_ex(id ID, extra_window_flags WindowFlags) bool

@[c: 'igBeginPopupMenuEx']
fn begin_popup_menu_ex(id ID, label &i8, extra_window_flags WindowFlags) bool

@[c: 'igOpenPopupEx']
fn open_popup_ex(id ID, popup_flags PopupFlags)

@[c: 'igClosePopupToLevel']
fn close_popup_to_level(remaining int, restore_focus_to_window_under_popup bool)

@[c: 'igClosePopupsOverWindow']
fn close_popups_over_window(ref_window &Window, restore_focus_to_window_under_popup bool)

@[c: 'igClosePopupsExceptModals']
fn close_popups_except_modals()

@[c: 'igIsPopupOpen_ID']
fn is_popup_open_id(id ID, popup_flags PopupFlags) bool

@[c: 'igGetPopupAllowedExtentRect']
fn get_popup_allowed_extent_rect(p_out &C.ImRect, window &Window)

@[c: 'igGetTopMostPopupModal']
fn get_top_most_popup_modal() &Window

@[c: 'igGetTopMostAndVisiblePopupModal']
fn get_top_most_and_visible_popup_modal() &Window

@[c: 'igFindBlockingModal']
fn find_blocking_modal(window &Window) &Window

@[c: 'igFindBestWindowPosForPopup']
fn find_best_window_pos_for_popup(p_out &ImVec2, window &Window)

@[c: 'igFindBestWindowPosForPopupEx']
fn find_best_window_pos_for_popup_ex(p_out &ImVec2, ref_pos ImVec2, size ImVec2, last_dir &Dir, r_outer C.ImRect, r_avoid C.ImRect, policy PopupPositionPolicy)

@[c: 'igBeginTooltipEx']
fn begin_tooltip_ex(tooltip_flags TooltipFlags, extra_window_flags WindowFlags) bool

@[c: 'igBeginTooltipHidden']
fn begin_tooltip_hidden() bool

@[c: 'igBeginViewportSideBar']
fn begin_viewport_side_bar(name &i8, viewport &Viewport, dir Dir, size f32, window_flags WindowFlags) bool

@[c: 'igBeginMenuEx']
fn begin_menu_ex(label &i8, icon &i8, enabled bool) bool

@[c: 'igMenuItemEx']
fn menu_item_ex(label &i8, icon &i8, shortcut &i8, selected bool, enabled bool) bool

@[c: 'igBeginComboPopup']
fn begin_combo_popup(popup_id ID, bb C.ImRect, flags ComboFlags) bool

@[c: 'igBeginComboPreview']
fn begin_combo_preview() bool

@[c: 'igEndComboPreview']
fn end_combo_preview()

@[c: 'igNavInitWindow']
fn nav_init_window(window &Window, force_reinit bool)

@[c: 'igNavInitRequestApplyResult']
fn nav_init_request_apply_result()

@[c: 'igNavMoveRequestButNoResultYet']
fn nav_move_request_but_no_result_yet() bool

@[c: 'igNavMoveRequestSubmit']
fn nav_move_request_submit(move_dir Dir, clip_dir Dir, move_flags NavMoveFlags, scroll_flags ScrollFlags)

@[c: 'igNavMoveRequestForward']
fn nav_move_request_forward(move_dir Dir, clip_dir Dir, move_flags NavMoveFlags, scroll_flags ScrollFlags)

@[c: 'igNavMoveRequestResolveWithLastItem']
fn nav_move_request_resolve_with_last_item(result &NavItemData)

@[c: 'igNavMoveRequestResolveWithPastTreeNode']
fn nav_move_request_resolve_with_past_tree_node(result &NavItemData, tree_node_data &TreeNodeStackData)

@[c: 'igNavMoveRequestCancel']
fn nav_move_request_cancel()

@[c: 'igNavMoveRequestApplyResult']
fn nav_move_request_apply_result()

@[c: 'igNavMoveRequestTryWrapping']
fn nav_move_request_try_wrapping(window &Window, move_flags NavMoveFlags)

@[c: 'igNavHighlightActivated']
fn nav_highlight_activated(id ID)

@[c: 'igNavClearPreferredPosForAxis']
fn nav_clear_preferred_pos_for_axis(axis Axis)

@[c: 'igSetNavCursorVisibleAfterMove']
fn set_nav_cursor_visible_after_move()

@[c: 'igNavUpdateCurrentWindowIsScrollPushableX']
fn nav_update_current_window_is_scroll_pushable_x()

@[c: 'igSetNavWindow']
fn set_nav_window(window &Window)

@[c: 'igSetNavID']
fn set_nav_id(id ID, nav_layer NavLayer, focus_scope_id ID, rect_rel C.ImRect)

@[c: 'igSetNavFocusScope']
fn set_nav_focus_scope(focus_scope_id ID)

@[c: 'igFocusItem']
fn focus_item()

@[c: 'igActivateItemByID']
fn activate_item_by_id(id ID)

@[c: 'igIsNamedKey']
fn is_named_key(key Key) bool

@[c: 'igIsNamedKeyOrMod']
fn is_named_key_or_mod(key Key) bool

@[c: 'igIsLegacyKey']
fn is_legacy_key(key Key) bool

@[c: 'igIsKeyboardKey']
fn is_keyboard_key(key Key) bool

@[c: 'igIsGamepadKey']
fn is_gamepad_key(key Key) bool

@[c: 'igIsMouseKey']
fn is_mouse_key(key Key) bool

@[c: 'igIsAliasKey']
fn is_alias_key(key Key) bool

@[c: 'igIsLRModKey']
fn is_lrm_od_key(key Key) bool

@[c: 'igFixupKeyChord']
fn fixup_key_chord(key_chord KeyChord) KeyChord

@[c: 'igConvertSingleModFlagToKey']
fn convert_single_mod_flag_to_key(key Key) Key

@[c: 'igGetKeyData_ContextPtr']
fn get_key_data_context_ptr(ctx &Context, key Key) &KeyData

@[c: 'igGetKeyData_Key']
fn get_key_data_key(key Key) &KeyData

@[c: 'igGetKeyChordName']
fn get_key_chord_name(key_chord KeyChord) &i8

@[c: 'igMouseButtonToKey']
fn mouse_button_to_key(button MouseButton) Key

@[c: 'igIsMouseDragPastThreshold']
fn is_mouse_drag_past_threshold(button MouseButton, lock_threshold f32) bool

@[c: 'igGetKeyMagnitude2d']
fn get_key_magnitude2d(p_out &ImVec2, key_left Key, key_right Key, key_up Key, key_down Key)

@[c: 'igGetNavTweakPressedAmount']
fn get_nav_tweak_pressed_amount(axis Axis) f32

@[c: 'igCalcTypematicRepeatAmount']
fn calc_typematic_repeat_amount(t0 f32, t1 f32, repeat_delay f32, repeat_rate f32) int

@[c: 'igGetTypematicRepeatRate']
fn get_typematic_repeat_rate(flags InputFlags, repeat_delay &f32, repeat_rate &f32)

@[c: 'igTeleportMousePos']
fn teleport_mouse_pos(pos ImVec2)

@[c: 'igSetActiveIdUsingAllKeyboardKeys']
fn set_active_id_using_all_keyboard_keys()

@[c: 'igIsActiveIdUsingNavDir']
fn is_active_id_using_nav_dir(dir Dir) bool

@[c: 'igGetKeyOwner']
fn get_key_owner(key Key) ID

@[c: 'igSetKeyOwner']
fn set_key_owner(key Key, owner_id ID, flags InputFlags)

@[c: 'igSetKeyOwnersForKeyChord']
fn set_key_owners_for_key_chord(key KeyChord, owner_id ID, flags InputFlags)

@[c: 'igSetItemKeyOwner_InputFlags']
fn set_item_key_owner_input_flags(key Key, flags InputFlags)

@[c: 'igTestKeyOwner']
fn test_key_owner(key Key, owner_id ID) bool

@[c: 'igGetKeyOwnerData']
fn get_key_owner_data(ctx &Context, key Key) &KeyOwnerData

@[c: 'igIsKeyDown_ID']
fn is_key_down_id(key Key, owner_id ID) bool

@[c: 'igIsKeyPressed_InputFlags']
fn is_key_pressed_input_flags(key Key, flags InputFlags, owner_id ID) bool

@[c: 'igIsKeyReleased_ID']
fn is_key_released_id(key Key, owner_id ID) bool

@[c: 'igIsKeyChordPressed_InputFlags']
fn is_key_chord_pressed_input_flags(key_chord KeyChord, flags InputFlags, owner_id ID) bool

@[c: 'igIsMouseDown_ID']
fn is_mouse_down_id(button MouseButton, owner_id ID) bool

@[c: 'igIsMouseClicked_InputFlags']
fn is_mouse_clicked_input_flags(button MouseButton, flags InputFlags, owner_id ID) bool

@[c: 'igIsMouseReleased_ID']
fn is_mouse_released_id(button MouseButton, owner_id ID) bool

@[c: 'igIsMouseDoubleClicked_ID']
fn is_mouse_double_clicked_id(button MouseButton, owner_id ID) bool

@[c: 'igShortcut_ID']
fn shortcut_id(key_chord KeyChord, flags InputFlags, owner_id ID) bool

@[c: 'igSetShortcutRouting']
fn set_shortcut_routing(key_chord KeyChord, flags InputFlags, owner_id ID) bool

@[c: 'igTestShortcutRouting']
fn test_shortcut_routing(key_chord KeyChord, owner_id ID) bool

@[c: 'igGetShortcutRoutingData']
fn get_shortcut_routing_data(key_chord KeyChord) &KeyRoutingData

@[c: 'igDockContextInitialize']
fn dock_context_initialize(ctx &Context)

@[c: 'igDockContextShutdown']
fn dock_context_shutdown(ctx &Context)

@[c: 'igDockContextClearNodes']
fn dock_context_clear_nodes(ctx &Context, root_id ID, clear_settings_refs bool)

@[c: 'igDockContextRebuildNodes']
fn dock_context_rebuild_nodes(ctx &Context)

@[c: 'igDockContextNewFrameUpdateUndocking']
fn dock_context_new_frame_update_undocking(ctx &Context)

@[c: 'igDockContextNewFrameUpdateDocking']
fn dock_context_new_frame_update_docking(ctx &Context)

@[c: 'igDockContextEndFrame']
fn dock_context_end_frame(ctx &Context)

@[c: 'igDockContextGenNodeID']
fn dock_context_gen_node_id(ctx &Context) ID

@[c: 'igDockContextQueueDock']
fn dock_context_queue_dock(ctx &Context, target &Window, target_node &DockNode, payload &Window, split_dir Dir, split_ratio f32, split_outer bool)

@[c: 'igDockContextQueueUndockWindow']
fn dock_context_queue_undock_window(ctx &Context, window &Window)

@[c: 'igDockContextQueueUndockNode']
fn dock_context_queue_undock_node(ctx &Context, node &DockNode)

@[c: 'igDockContextProcessUndockWindow']
fn dock_context_process_undock_window(ctx &Context, window &Window, clear_persistent_docking_ref bool)

@[c: 'igDockContextProcessUndockNode']
fn dock_context_process_undock_node(ctx &Context, node &DockNode)

@[c: 'igDockContextCalcDropPosForDocking']
fn dock_context_calc_drop_pos_for_docking(target &Window, target_node &DockNode, payload_window &Window, payload_node &DockNode, split_dir Dir, split_outer bool, out_pos &ImVec2) bool

@[c: 'igDockContextFindNodeByID']
fn dock_context_find_node_by_id(ctx &Context, id ID) &DockNode

@[c: 'igDockNodeWindowMenuHandler_Default']
fn dock_node_window_menu_handler_default(ctx &Context, node &DockNode, tab_bar &C.ImGuiTabBar)

@[c: 'igDockNodeBeginAmendTabBar']
fn dock_node_begin_amend_tab_bar(node &DockNode) bool

@[c: 'igDockNodeEndAmendTabBar']
fn dock_node_end_amend_tab_bar()

@[c: 'igDockNodeGetRootNode']
fn dock_node_get_root_node(node &DockNode) &DockNode

@[c: 'igDockNodeIsInHierarchyOf']
fn dock_node_is_in_hierarchy_of(node &DockNode, parent &DockNode) bool

@[c: 'igDockNodeGetDepth']
fn dock_node_get_depth(node &DockNode) int

@[c: 'igDockNodeGetWindowMenuButtonId']
fn dock_node_get_window_menu_button_id(node &DockNode) ID

@[c: 'igGetWindowDockNode']
fn get_window_dock_node() &DockNode

@[c: 'igGetWindowAlwaysWantOwnTabBar']
fn get_window_always_want_own_tab_bar(window &Window) bool

@[c: 'igBeginDocked']
fn begin_docked(window &Window, p_open &bool)

@[c: 'igBeginDockableDragDropSource']
fn begin_dockable_drag_drop_source(window &Window)

@[c: 'igBeginDockableDragDropTarget']
fn begin_dockable_drag_drop_target(window &Window)

@[c: 'igSetWindowDock']
fn set_window_dock(window &Window, dock_id ID, cond Cond)

@[c: 'igDockBuilderDockWindow']
fn dock_builder_dock_window(window_name &i8, node_id ID)

@[c: 'igDockBuilderGetNode']
fn dock_builder_get_node(node_id ID) &DockNode

@[c: 'igDockBuilderGetCentralNode']
fn dock_builder_get_central_node(node_id ID) &DockNode

@[c: 'igDockBuilderAddNode']
fn dock_builder_add_node(node_id ID, flags DockNodeFlags) ID

@[c: 'igDockBuilderRemoveNode']
fn dock_builder_remove_node(node_id ID)

@[c: 'igDockBuilderRemoveNodeDockedWindows']
fn dock_builder_remove_node_docked_windows(node_id ID, clear_settings_refs bool)

@[c: 'igDockBuilderRemoveNodeChildNodes']
fn dock_builder_remove_node_child_nodes(node_id ID)

@[c: 'igDockBuilderSetNodePos']
fn dock_builder_set_node_pos(node_id ID, pos ImVec2)

@[c: 'igDockBuilderSetNodeSize']
fn dock_builder_set_node_size(node_id ID, size ImVec2)

@[c: 'igDockBuilderSplitNode']
fn dock_builder_split_node(node_id ID, split_dir Dir, size_ratio_for_node_at_dir f32, out_id_at_dir &ID, out_id_at_opposite_dir &ID) ID

@[c: 'igDockBuilderCopyDockSpace']
fn dock_builder_copy_dock_space(src_dockspace_id ID, dst_dockspace_id ID, in_window_remap_pairs &ImVector_const_charPtr)

@[c: 'igDockBuilderCopyNode']
fn dock_builder_copy_node(src_node_id ID, dst_node_id ID, out_node_remap_pairs &ImVector_ImGuiID)

@[c: 'igDockBuilderCopyWindowSettings']
fn dock_builder_copy_window_settings(src_name &i8, dst_name &i8)

@[c: 'igDockBuilderFinish']
fn dock_builder_finish(node_id ID)

@[c: 'igPushFocusScope']
fn push_focus_scope(id ID)

@[c: 'igPopFocusScope']
fn pop_focus_scope()

@[c: 'igGetCurrentFocusScope']
fn get_current_focus_scope() ID

@[c: 'igIsDragDropActive']
fn is_drag_drop_active() bool

@[c: 'igBeginDragDropTargetCustom']
fn begin_drag_drop_target_custom(bb C.ImRect, id ID) bool

@[c: 'igClearDragDrop']
fn clear_drag_drop()

@[c: 'igIsDragDropPayloadBeingAccepted']
fn is_drag_drop_payload_being_accepted() bool

@[c: 'igRenderDragDropTargetRect']
fn render_drag_drop_target_rect(bb C.ImRect, item_clip_rect C.ImRect)

@[c: 'igGetTypingSelectRequest']
fn get_typing_select_request(flags TypingSelectFlags) &TypingSelectRequest

@[c: 'igTypingSelectFindMatch']
fn typing_select_find_match(req &TypingSelectRequest, items_count int, get_item_name_func fn (voidptr, int) &i8, user_data voidptr, nav_item_idx int) int

@[c: 'igTypingSelectFindNextSingleCharMatch']
fn typing_select_find_next_single_char_match(req &TypingSelectRequest, items_count int, get_item_name_func fn (voidptr, int) &i8, user_data voidptr, nav_item_idx int) int

@[c: 'igTypingSelectFindBestLeadingMatch']
fn typing_select_find_best_leading_match(req &TypingSelectRequest, items_count int, get_item_name_func fn (voidptr, int) &i8, user_data voidptr) int

@[c: 'igBeginBoxSelect']
fn begin_box_select(scope_rect C.ImRect, window &Window, box_select_id ID, ms_flags MultiSelectFlags) bool

@[c: 'igEndBoxSelect']
fn end_box_select(scope_rect C.ImRect, ms_flags MultiSelectFlags)

@[c: 'igMultiSelectItemHeader']
fn multi_select_item_header(id ID, p_selected &bool, p_button_flags &ButtonFlags)

@[c: 'igMultiSelectItemFooter']
fn multi_select_item_footer(id ID, p_selected &bool, p_pressed &bool)

@[c: 'igMultiSelectAddSetAll']
fn multi_select_add_set_all(ms &MultiSelectTempData, selected bool)

@[c: 'igMultiSelectAddSetRange']
fn multi_select_add_set_range(ms &MultiSelectTempData, selected bool, range_dir int, first_item SelectionUserData, last_item SelectionUserData)

@[c: 'igGetBoxSelectState']
fn get_box_select_state(id ID) &BoxSelectState

@[c: 'igGetMultiSelectState']
fn get_multi_select_state(id ID) &MultiSelectState

@[c: 'igSetWindowClipRectBeforeSetChannel']
fn set_window_clip_rect_before_set_channel(window &Window, clip_rect C.ImRect)

@[c: 'igBeginColumns']
fn begin_columns(str_id &i8, count int, flags OldColumnFlags)

@[c: 'igEndColumns']
fn end_columns()

@[c: 'igPushColumnClipRect']
fn push_column_clip_rect(column_index int)

@[c: 'igPushColumnsBackground']
fn push_columns_background()

@[c: 'igPopColumnsBackground']
fn pop_columns_background()

@[c: 'igGetColumnsID']
fn get_columns_id(str_id &i8, count int) ID

@[c: 'igFindOrCreateColumns']
fn find_or_create_columns(window &Window, id ID) &OldColumns

@[c: 'igGetColumnOffsetFromNorm']
fn get_column_offset_from_norm(columns &OldColumns, offset_norm f32) f32

@[c: 'igGetColumnNormFromOffset']
fn get_column_norm_from_offset(columns &OldColumns, offset f32) f32

@[c: 'igTableOpenContextMenu']
fn table_open_context_menu(column_n int)

@[c: 'igTableSetColumnWidth']
fn table_set_column_width(column_n int, width f32)

@[c: 'igTableSetColumnSortDirection']
fn table_set_column_sort_direction(column_n int, sort_direction SortDirection, append_to_sort_specs bool)

@[c: 'igTableGetHoveredRow']
fn table_get_hovered_row() int

@[c: 'igTableGetHeaderRowHeight']
fn table_get_header_row_height() f32

@[c: 'igTableGetHeaderAngledMaxLabelWidth']
fn table_get_header_angled_max_label_width() f32

@[c: 'igTablePushBackgroundChannel']
fn table_push_background_channel()

@[c: 'igTablePopBackgroundChannel']
fn table_pop_background_channel()

@[c: 'igTableAngledHeadersRowEx']
fn table_angled_headers_row_ex(row_id ID, angle f32, max_label_width f32, data &TableHeaderData, data_count int)

@[c: 'igGetCurrentTable']
fn get_current_table() &Table

@[c: 'igTableFindByID']
fn table_find_by_id(id ID) &Table

@[c: 'igBeginTableEx']
fn begin_table_ex(name &i8, id ID, columns_count int, flags TableFlags, outer_size ImVec2, inner_width f32) bool

@[c: 'igTableBeginInitMemory']
fn table_begin_init_memory(table &Table, columns_count int)

@[c: 'igTableBeginApplyRequests']
fn table_begin_apply_requests(table &Table)

@[c: 'igTableSetupDrawChannels']
fn table_setup_draw_channels(table &Table)

@[c: 'igTableUpdateLayout']
fn table_update_layout(table &Table)

@[c: 'igTableUpdateBorders']
fn table_update_borders(table &Table)

@[c: 'igTableUpdateColumnsWeightFromWidth']
fn table_update_columns_weight_from_width(table &Table)

@[c: 'igTableDrawBorders']
fn table_draw_borders(table &Table)

@[c: 'igTableDrawDefaultContextMenu']
fn table_draw_default_context_menu(table &Table, flags_for_section_to_display TableFlags)

@[c: 'igTableBeginContextMenuPopup']
fn table_begin_context_menu_popup(table &Table) bool

@[c: 'igTableMergeDrawChannels']
fn table_merge_draw_channels(table &Table)

@[c: 'igTableGetInstanceData']
fn table_get_instance_data(table &Table, instance_no int) &TableInstanceData

@[c: 'igTableGetInstanceID']
fn table_get_instance_id(table &Table, instance_no int) ID

@[c: 'igTableSortSpecsSanitize']
fn table_sort_specs_sanitize(table &Table)

@[c: 'igTableSortSpecsBuild']
fn table_sort_specs_build(table &Table)

@[c: 'igTableGetColumnNextSortDirection']
fn table_get_column_next_sort_direction(column &TableColumn) SortDirection

@[c: 'igTableFixColumnSortDirection']
fn table_fix_column_sort_direction(table &Table, column &TableColumn)

@[c: 'igTableGetColumnWidthAuto']
fn table_get_column_width_auto(table &Table, column &TableColumn) f32

@[c: 'igTableBeginRow']
fn table_begin_row(table &Table)

@[c: 'igTableEndRow']
fn table_end_row(table &Table)

@[c: 'igTableBeginCell']
fn table_begin_cell(table &Table, column_n int)

@[c: 'igTableEndCell']
fn table_end_cell(table &Table)

@[c: 'igTableGetCellBgRect']
fn table_get_cell_bg_rect(p_out &C.ImRect, table &Table, column_n int)

@[c: 'igTableGetColumnName_TablePtr']
fn table_get_column_name_table_ptr(table &Table, column_n int) &i8

@[c: 'igTableGetColumnResizeID']
fn table_get_column_resize_id(table &Table, column_n int, instance_no int) ID

@[c: 'igTableCalcMaxColumnWidth']
fn table_calc_max_column_width(table &Table, column_n int) f32

@[c: 'igTableSetColumnWidthAutoSingle']
fn table_set_column_width_auto_single(table &Table, column_n int)

@[c: 'igTableSetColumnWidthAutoAll']
fn table_set_column_width_auto_all(table &Table)

@[c: 'igTableRemove']
fn table_remove(table &Table)

@[c: 'igTableGcCompactTransientBuffers_TablePtr']
fn table_gc_compact_transient_buffers_table_ptr(table &Table)

@[c: 'igTableGcCompactTransientBuffers_TableTempDataPtr']
fn table_gc_compact_transient_buffers_table_temp_data_ptr(table &TableTempData)

@[c: 'igTableGcCompactSettings']
fn table_gc_compact_settings()

@[c: 'igTableLoadSettings']
fn table_load_settings(table &Table)

@[c: 'igTableSaveSettings']
fn table_save_settings(table &Table)

@[c: 'igTableResetSettings']
fn table_reset_settings(table &Table)

@[c: 'igTableGetBoundSettings']
fn table_get_bound_settings(table &Table) &TableSettings

@[c: 'igTableSettingsAddSettingsHandler']
fn table_settings_add_settings_handler()

@[c: 'igTableSettingsCreate']
fn table_settings_create(id ID, columns_count int) &TableSettings

@[c: 'igTableSettingsFindByID']
fn table_settings_find_by_id(id ID) &TableSettings

@[c: 'igGetCurrentTabBar']
fn get_current_tab_bar() &C.ImGuiTabBar

@[c: 'igBeginTabBarEx']
fn begin_tab_bar_ex(tab_bar &C.ImGuiTabBar, bb C.ImRect, flags ImGuiTabBarFlags) bool

@[c: 'igTabBarFindTabByID']
fn tab_bar_find_tab_by_id(tab_bar &C.ImGuiTabBar, tab_id ID) &TabItem

@[c: 'igTabBarFindTabByOrder']
fn tab_bar_find_tab_by_order(tab_bar &C.ImGuiTabBar, order int) &TabItem

@[c: 'igTabBarFindMostRecentlySelectedTabForActiveWindow']
fn tab_bar_find_most_recently_selected_tab_for_active_window(tab_bar &C.ImGuiTabBar) &TabItem

@[c: 'igTabBarGetCurrentTab']
fn tab_bar_get_current_tab(tab_bar &C.ImGuiTabBar) &TabItem

@[c: 'igTabBarGetTabOrder']
fn tab_bar_get_tab_order(tab_bar &C.ImGuiTabBar, tab &TabItem) int

@[c: 'igTabBarGetTabName']
fn tab_bar_get_tab_name(tab_bar &C.ImGuiTabBar, tab &TabItem) &i8

@[c: 'igTabBarAddTab']
fn tab_bar_add_tab(tab_bar &C.ImGuiTabBar, tab_flags TabItemFlags, window &Window)

@[c: 'igTabBarRemoveTab']
fn tab_bar_remove_tab(tab_bar &C.ImGuiTabBar, tab_id ID)

@[c: 'igTabBarCloseTab']
fn tab_bar_close_tab(tab_bar &C.ImGuiTabBar, tab &TabItem)

@[c: 'igTabBarQueueFocus_TabItemPtr']
fn tab_bar_queue_focus_tab_item_ptr(tab_bar &C.ImGuiTabBar, tab &TabItem)

@[c: 'igTabBarQueueFocus_Str']
fn tab_bar_queue_focus_str(tab_bar &C.ImGuiTabBar, tab_name &i8)

@[c: 'igTabBarQueueReorder']
fn tab_bar_queue_reorder(tab_bar &C.ImGuiTabBar, tab &TabItem, offset int)

@[c: 'igTabBarQueueReorderFromMousePos']
fn tab_bar_queue_reorder_from_mouse_pos(tab_bar &C.ImGuiTabBar, tab &TabItem, mouse_pos ImVec2)

@[c: 'igTabBarProcessReorder']
fn tab_bar_process_reorder(tab_bar &C.ImGuiTabBar) bool

@[c: 'igTabItemEx']
fn tab_item_ex(tab_bar &C.ImGuiTabBar, label &i8, p_open &bool, flags TabItemFlags, docked_window &Window) bool

@[c: 'igTabItemSpacing']
fn tab_item_spacing(str_id &i8, flags TabItemFlags, width f32)

@[c: 'igTabItemCalcSize_Str']
fn tab_item_calc_size_str(p_out &ImVec2, label &i8, has_close_button_or_unsaved_marker bool)

@[c: 'igTabItemCalcSize_WindowPtr']
fn tab_item_calc_size_window_ptr(p_out &ImVec2, window &Window)

@[c: 'igTabItemBackground']
fn tab_item_background(draw_list &ImDrawList, bb C.ImRect, flags TabItemFlags, col ImU32)

@[c: 'igTabItemLabelAndCloseButton']
fn tab_item_label_and_close_button(draw_list &ImDrawList, bb C.ImRect, flags TabItemFlags, frame_padding ImVec2, label &i8, tab_id ID, close_button_id ID, is_contents_visible bool, out_just_closed &bool, out_text_clipped &bool)

@[c: 'igRenderText']
fn render_text(pos ImVec2, text &i8, text_end &i8, hide_text_after_hash bool)

@[c: 'igRenderTextWrapped']
fn render_text_wrapped(pos ImVec2, text &i8, text_end &i8, wrap_width f32)

@[c: 'igRenderTextClipped']
fn render_text_clipped(pos_min ImVec2, pos_max ImVec2, text &i8, text_end &i8, text_size_if_known &ImVec2, align ImVec2, clip_rect &C.ImRect)

@[c: 'igRenderTextClippedEx']
fn render_text_clipped_ex(draw_list &ImDrawList, pos_min ImVec2, pos_max ImVec2, text &i8, text_end &i8, text_size_if_known &ImVec2, align ImVec2, clip_rect &C.ImRect)

@[c: 'igRenderTextEllipsis']
fn render_text_ellipsis(draw_list &ImDrawList, pos_min ImVec2, pos_max ImVec2, clip_max_x f32, ellipsis_max_x f32, text &i8, text_end &i8, text_size_if_known &ImVec2)

@[c: 'igRenderFrame']
fn render_frame(p_min ImVec2, p_max ImVec2, fill_col ImU32, borders bool, rounding f32)

@[c: 'igRenderFrameBorder']
fn render_frame_border(p_min ImVec2, p_max ImVec2, rounding f32)

@[c: 'igRenderColorRectWithAlphaCheckerboard']
fn render_color_rect_with_alpha_checkerboard(draw_list &ImDrawList, p_min ImVec2, p_max ImVec2, fill_col ImU32, grid_step f32, grid_off ImVec2, rounding f32, flags ImDrawFlags)

@[c: 'igRenderNavCursor']
fn render_nav_cursor(bb C.ImRect, id ID, flags NavRenderCursorFlags)

@[c: 'igFindRenderedTextEnd']
fn find_rendered_text_end(text &i8, text_end &i8) &i8

@[c: 'igRenderMouseCursor']
fn render_mouse_cursor(pos ImVec2, scale f32, mouse_cursor MouseCursor, col_fill ImU32, col_border ImU32, col_shadow ImU32)

@[c: 'igRenderArrow']
fn render_arrow(draw_list &ImDrawList, pos ImVec2, col ImU32, dir Dir, scale f32)

@[c: 'igRenderBullet']
fn render_bullet(draw_list &ImDrawList, pos ImVec2, col ImU32)

@[c: 'igRenderCheckMark']
fn render_check_mark(draw_list &ImDrawList, pos ImVec2, col ImU32, sz f32)

@[c: 'igRenderArrowPointingAt']
fn render_arrow_pointing_at(draw_list &ImDrawList, pos ImVec2, half_sz ImVec2, direction Dir, col ImU32)

@[c: 'igRenderArrowDockMenu']
fn render_arrow_dock_menu(draw_list &ImDrawList, p_min ImVec2, sz f32, col ImU32)

@[c: 'igRenderRectFilledRangeH']
fn render_rect_filled_range_h(draw_list &ImDrawList, rect C.ImRect, col ImU32, x_start_norm f32, x_end_norm f32, rounding f32)

@[c: 'igRenderRectFilledWithHole']
fn render_rect_filled_with_hole(draw_list &ImDrawList, outer C.ImRect, inner C.ImRect, col ImU32, rounding f32)

@[c: 'igCalcRoundingFlagsForRectInRect']
fn calc_rounding_flags_for_rect_in_rect(r_in C.ImRect, r_outer C.ImRect, threshold f32) ImDrawFlags

@[c: 'igTextEx']
fn text_ex(text &i8, text_end &i8, flags TextFlags)

@[c: 'igButtonEx']
fn button_ex(label &i8, size_arg ImVec2, flags ButtonFlags) bool

@[c: 'igArrowButtonEx']
fn arrow_button_ex(str_id &i8, dir Dir, size_arg ImVec2, flags ButtonFlags) bool

@[c: 'igImageButtonEx']
fn image_button_ex(id ID, user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col C.ImVec4, tint_col C.ImVec4, flags ButtonFlags) bool

@[c: 'igSeparatorEx']
fn separator_ex(flags SeparatorFlags, thickness f32)

@[c: 'igSeparatorTextEx']
fn separator_text_ex(id ID, label &i8, label_end &i8, extra_width f32)

@[c: 'igCheckboxFlags_S64Ptr']
fn checkbox_flags_s64_ptr(label &i8, flags &ImS64, flags_value ImS64) bool

@[c: 'igCheckboxFlags_U64Ptr']
fn checkbox_flags_u64_ptr(label &i8, flags &ImU64, flags_value ImU64) bool

@[c: 'igCloseButton']
fn close_button(id ID, pos ImVec2) bool

@[c: 'igCollapseButton']
fn collapse_button(id ID, pos ImVec2, dock_node &DockNode) bool

@[c: 'igScrollbar']
fn scrollbar(axis Axis)

@[c: 'igScrollbarEx']
fn scrollbar_ex(bb C.ImRect, id ID, axis Axis, p_scroll_v &ImS64, avail_v ImS64, contents_v ImS64, draw_rounding_flags ImDrawFlags) bool

@[c: 'igGetWindowScrollbarRect']
fn get_window_scrollbar_rect(p_out &C.ImRect, window &Window, axis Axis)

@[c: 'igGetWindowScrollbarID']
fn get_window_scrollbar_id(window &Window, axis Axis) ID

@[c: 'igGetWindowResizeCornerID']
fn get_window_resize_corner_id(window &Window, n int) ID

@[c: 'igGetWindowResizeBorderID']
fn get_window_resize_border_id(window &Window, dir Dir) ID

@[c: 'igButtonBehavior']
fn button_behavior(bb C.ImRect, id ID, out_hovered &bool, out_held &bool, flags ButtonFlags) bool

@[c: 'igDragBehavior']
fn drag_behavior(id ID, data_type DataType, p_v voidptr, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igSliderBehavior']
fn slider_behavior(bb C.ImRect, id ID, data_type DataType, p_v voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags, out_grab_bb &C.ImRect) bool

@[c: 'igSplitterBehavior']
fn splitter_behavior(bb C.ImRect, id ID, axis Axis, size1 &f32, size2 &f32, min_size1 f32, min_size2 f32, hover_extend f32, hover_visibility_delay f32, bg_col ImU32) bool

@[c: 'igTreeNodeBehavior']
fn tree_node_behavior(id ID, flags TreeNodeFlags, label &i8, label_end &i8) bool

@[c: 'igTreePushOverrideID']
fn tree_push_override_id(id ID)

@[c: 'igTreeNodeGetOpen']
fn tree_node_get_open(storage_id ID) bool

@[c: 'igTreeNodeSetOpen']
fn tree_node_set_open(storage_id ID, open bool)

@[c: 'igTreeNodeUpdateNextOpen']
fn tree_node_update_next_open(storage_id ID, flags TreeNodeFlags) bool

@[c: 'igDataTypeGetInfo']
fn data_type_get_info(data_type DataType) &DataTypeInfo

@[c: 'igDataTypeFormatString']
fn data_type_format_string(buf &i8, buf_size int, data_type DataType, p_data voidptr, format &i8) int

@[c: 'igDataTypeApplyOp']
fn data_type_apply_op(data_type DataType, op int, output voidptr, arg_1 voidptr, arg_2 voidptr)

@[c: 'igDataTypeApplyFromText']
fn data_type_apply_from_text(buf &i8, data_type DataType, p_data voidptr, format &i8, p_data_when_empty voidptr) bool

@[c: 'igDataTypeCompare']
fn data_type_compare(data_type DataType, arg_1 voidptr, arg_2 voidptr) int

@[c: 'igDataTypeClamp']
fn data_type_clamp(data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr) bool

@[c: 'igDataTypeIsZero']
fn data_type_is_zero(data_type DataType, p_data voidptr) bool

@[c: 'igInputTextEx']
fn input_text_ex(label &i8, hint &i8, buf &i8, buf_size int, size_arg ImVec2, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c: 'igInputTextDeactivateHook']
fn input_text_deactivate_hook(id ID)

@[c: 'igTempInputText']
fn temp_input_text(bb C.ImRect, id ID, label &i8, buf &i8, buf_size int, flags InputTextFlags) bool

@[c: 'igTempInputScalar']
fn temp_input_scalar(bb C.ImRect, id ID, label &i8, data_type DataType, p_data voidptr, format &i8, p_clamp_min voidptr, p_clamp_max voidptr) bool

@[c: 'igTempInputIsActive']
fn temp_input_is_active(id ID) bool

@[c: 'igGetInputTextState']
fn get_input_text_state(id ID) &InputTextState

@[c: 'igSetNextItemRefVal']
fn set_next_item_ref_val(data_type DataType, p_data voidptr)

@[c: 'igIsItemActiveAsInputText']
fn is_item_active_as_input_text() bool

@[c: 'igColorTooltip']
fn color_tooltip(text &i8, col &f32, flags ColorEditFlags)

@[c: 'igColorEditOptionsPopup']
fn color_edit_options_popup(col &f32, flags ColorEditFlags)

@[c: 'igColorPickerOptionsPopup']
fn color_picker_options_popup(ref_col &f32, flags ColorEditFlags)

@[c: 'igPlotEx']
fn plot_ex(plot_type PlotType, label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, size_arg ImVec2) int

@[c: 'igShadeVertsLinearColorGradientKeepAlpha']
fn shade_verts_linear_color_gradient_keep_alpha(draw_list &ImDrawList, vert_start_idx int, vert_end_idx int, gradient_p0 ImVec2, gradient_p1 ImVec2, col0 ImU32, col1 ImU32)

@[c: 'igShadeVertsLinearUV']
fn shade_verts_linear_uv(draw_list &ImDrawList, vert_start_idx int, vert_end_idx int, a ImVec2, b ImVec2, uv_a ImVec2, uv_b ImVec2, clamp bool)

@[c: 'igShadeVertsTransformPos']
fn shade_verts_transform_pos(draw_list &ImDrawList, vert_start_idx int, vert_end_idx int, pivot_in ImVec2, cos_a f32, sin_a f32, pivot_out ImVec2)

@[c: 'igGcCompactTransientMiscBuffers']
fn gc_compact_transient_misc_buffers()

@[c: 'igGcCompactTransientWindowBuffers']
fn gc_compact_transient_window_buffers(window &Window)

@[c: 'igGcAwakeTransientWindowBuffers']
fn gc_awake_transient_window_buffers(window &Window)

@[c: 'igErrorLog']
fn error_log(msg &i8) bool

@[c: 'igErrorRecoveryStoreState']
fn error_recovery_store_state(state_out &ErrorRecoveryState)

@[c: 'igErrorRecoveryTryToRecoverState']
fn error_recovery_try_to_recover_state(state_in &ErrorRecoveryState)

@[c: 'igErrorRecoveryTryToRecoverWindowState']
fn error_recovery_try_to_recover_window_state(state_in &ErrorRecoveryState)

@[c: 'igErrorCheckUsingSetCursorPosToExtendParentBoundaries']
fn error_check_using_set_cursor_pos_to_extend_parent_boundaries()

@[c: 'igErrorCheckEndFrameFinalizeErrorTooltip']
fn error_check_end_frame_finalize_error_tooltip()

@[c: 'igBeginErrorTooltip']
fn begin_error_tooltip() bool

@[c: 'igEndErrorTooltip']
fn end_error_tooltip()

@[c: 'igDebugAllocHook']
fn debug_alloc_hook(info &DebugAllocInfo, frame_count int, ptr voidptr, size usize)

@[c: 'igDebugDrawCursorPos']
fn debug_draw_cursor_pos(col ImU32)

@[c: 'igDebugDrawLineExtents']
fn debug_draw_line_extents(col ImU32)

@[c: 'igDebugDrawItemRect']
fn debug_draw_item_rect(col ImU32)

@[c: 'igDebugTextUnformattedWithLocateItem']
fn debug_text_unformatted_with_locate_item(line_begin &i8, line_end &i8)

@[c: 'igDebugLocateItem']
fn debug_locate_item(target_id ID)

@[c: 'igDebugLocateItemOnHover']
fn debug_locate_item_on_hover(target_id ID)

@[c: 'igDebugLocateItemResolveWithLastItem']
fn debug_locate_item_resolve_with_last_item()

@[c: 'igDebugBreakClearData']
fn debug_break_clear_data()

@[c: 'igDebugBreakButton']
fn debug_break_button(label &i8, description_of_location &i8) bool

@[c: 'igDebugBreakButtonTooltip']
fn debug_break_button_tooltip(keyboard_only bool, description_of_location &i8)

@[c: 'igShowFontAtlas']
fn show_font_atlas(atlas &ImFontAtlas)

@[c: 'igDebugHookIdInfo']
fn debug_hook_id_info(id ID, data_type DataType, data_id voidptr, data_id_end voidptr)

@[c: 'igDebugNodeColumns']
fn debug_node_columns(columns &OldColumns)

@[c: 'igDebugNodeDockNode']
fn debug_node_dock_node(node &DockNode, label &i8)

@[c: 'igDebugNodeDrawList']
fn debug_node_draw_list(window &Window, viewport &ViewportP, draw_list &ImDrawList, label &i8)

@[c: 'igDebugNodeDrawCmdShowMeshAndBoundingBox']
fn debug_node_draw_cmd_show_mesh_and_bounding_box(out_draw_list &ImDrawList, draw_list &ImDrawList, draw_cmd &ImDrawCmd, show_mesh bool, show_aabb bool)

@[c: 'igDebugNodeFont']
fn debug_node_font(font &ImFont)

@[c: 'igDebugNodeFontGlyph']
fn debug_node_font_glyph(font &ImFont, glyph &ImFontGlyph)

@[c: 'igDebugNodeStorage']
fn debug_node_storage(storage &Storage, label &i8)

@[c: 'igDebugNodeTabBar']
fn debug_node_tab_bar(tab_bar &C.ImGuiTabBar, label &i8)

@[c: 'igDebugNodeTable']
fn debug_node_table(table &Table)

@[c: 'igDebugNodeTableSettings']
fn debug_node_table_settings(settings &TableSettings)

@[c: 'igDebugNodeInputTextState']
fn debug_node_input_text_state(state &InputTextState)

@[c: 'igDebugNodeTypingSelectState']
fn debug_node_typing_select_state(state &TypingSelectState)

@[c: 'igDebugNodeMultiSelectState']
fn debug_node_multi_select_state(state &MultiSelectState)

@[c: 'igDebugNodeWindow']
fn debug_node_window(window &Window, label &i8)

@[c: 'igDebugNodeWindowSettings']
fn debug_node_window_settings(settings &WindowSettings)

@[c: 'igDebugNodeWindowsList']
fn debug_node_windows_list(windows &ImVector_ImGuiWindowPtr, label &i8)

@[c: 'igDebugNodeWindowsListByBeginStackParent']
fn debug_node_windows_list_by_begin_stack_parent(windows &&Window, windows_size int, parent_in_begin_stack &Window)

@[c: 'igDebugNodeViewport']
fn debug_node_viewport(viewport &ViewportP)

@[c: 'igDebugNodePlatformMonitor']
fn debug_node_platform_monitor(monitor &PlatformMonitor, label &i8, idx int)

@[c: 'igDebugRenderKeyboardPreview']
fn debug_render_keyboard_preview(draw_list &ImDrawList)

@[c: 'igDebugRenderViewportThumbnail']
fn debug_render_viewport_thumbnail(draw_list &ImDrawList, viewport &ViewportP, bb C.ImRect)

@[c: 'igImFontAtlasGetBuilderForStbTruetype']
fn im_font_atlas_get_builder_for_stb_truetype() &ImFontBuilderIO

@[c: 'igImFontAtlasUpdateSourcesPointers']
fn im_font_atlas_update_sources_pointers(atlas &ImFontAtlas)

@[c: 'igImFontAtlasBuildInit']
fn im_font_atlas_build_init(atlas &ImFontAtlas)

@[c: 'igImFontAtlasBuildSetupFont']
fn im_font_atlas_build_setup_font(atlas &ImFontAtlas, font &ImFont, src &ImFontConfig, ascent f32, descent f32)

@[c: 'igImFontAtlasBuildPackCustomRects']
fn im_font_atlas_build_pack_custom_rects(atlas &ImFontAtlas, stbrp_context_opaque voidptr)

@[c: 'igImFontAtlasBuildFinish']
fn im_font_atlas_build_finish(atlas &ImFontAtlas)

@[c: 'igImFontAtlasBuildRender8bppRectFromString']
fn im_font_atlas_build_render8bpp_rect_from_string(atlas &ImFontAtlas, x int, y int, w int, h int, in_str &i8, in_marker_char i8, in_marker_pixel_value u8)

@[c: 'igImFontAtlasBuildRender32bppRectFromString']
fn im_font_atlas_build_render32bpp_rect_from_string(atlas &ImFontAtlas, x int, y int, w int, h int, in_str &i8, in_marker_char i8, in_marker_pixel_value u32)

@[c: 'igImFontAtlasBuildMultiplyCalcLookupTable']
fn im_font_atlas_build_multiply_calc_lookup_table(out_table &u8, in_multiply_factor f32)

@[c: 'igImFontAtlasBuildMultiplyRectAlpha8']
fn im_font_atlas_build_multiply_rect_alpha8(table &u8, pixels &u8, x int, y int, w int, h int, stride int)

@[c: 'igImFontAtlasBuildGetOversampleFactors']
fn im_font_atlas_build_get_oversample_factors(src &ImFontConfig, out_oversample_h &int, out_oversample_v &int)

@[c: 'igImFontAtlasGetMouseCursorTexData']
fn im_font_atlas_get_mouse_cursor_tex_data(atlas &ImFontAtlas, cursor_type MouseCursor, out_offset &ImVec2, out_size &ImVec2, out_uv_border &ImVec2, out_uv_fill &ImVec2) bool

/////////////////////////hand written functions
// no LogTextV
@[c: 'igLogText']
@[c2v_variadic]
fn log_text(fmt ...&i8)

// no appendfV
@[c: 'ImGuiTextBuffer_appendf']
@[c2v_variadic]
fn text_buffer_appendf(self &TextBuffer, fmt ...&i8)

// for getting FLT_MAX in bindings
@[c: 'igGET_FLT_MAX']
fn get_flt_max() f32

// for getting FLT_MIN in bindings
@[c: 'igGET_FLT_MIN']
fn get_flt_min() f32

@[c: 'ImVector_ImWchar_create']
fn im_vector_im_wchar_create() &ImVector_ImWchar

@[c: 'ImVector_ImWchar_destroy']
fn im_vector_im_wchar_destroy(self &ImVector_ImWchar)

@[c: 'ImVector_ImWchar_Init']
fn im_vector_im_wchar_init(p &ImVector_ImWchar)

@[c: 'ImVector_ImWchar_UnInit']
fn im_vector_im_wchar_un_init(p &ImVector_ImWchar)

@[c: 'ImGuiPlatformIO_Set_Platform_GetWindowPos']
fn platform_io_set_platform_get_window_pos(platform_io &PlatformIO, user_callback fn (&Viewport, ImVec2))

@[c: 'ImGuiPlatformIO_Set_Platform_GetWindowSize']
fn platform_io_set_platform_get_window_size(platform_io &PlatformIO, user_callback fn (&Viewport, ImVec2))

// CIMGUI_INCLUDED
