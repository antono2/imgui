module implot
/*
#flag -I /home/anton/.vmodules/imgui/include

#include "time.h"

#include "cimplot.h"

#flag -DIMGUI_USE_WCHAR32
#flag -L /home/anton/.vmodules/imgui/lib
#flag -l cimplot
*/
