module imgui


#flag -I @VMODROOT/include
#flag -L @VMODROOT/lib
#flag -l :cimgui.a
#flag -l m
#flag -l stdc++

#define CIMGUI_DEFINE_ENUMS_AND_STRUCTS
#include "cimgui.h"

