/* 
  This contains things that were not automatically translated.
  Note that code is read by cleanup.perl and commented code is not ignored.
*/

module imgui
