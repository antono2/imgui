module imgui

#flag -l :cimplot.a

#include "time.h"
#include "cimplot.h"

