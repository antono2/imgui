module implot
/*
#flag -I @VMODROOT/include

#include "time.h"

#include "cimplot.h"

#flag -DIMGUI_USE_WCHAR32
#flag -L @VMODROOT/lib
#flag -Wl,-rpath=@VMODROOT/lib
#flag -l cimplot
*/
