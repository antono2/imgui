@[translated]
module imgui

#flag -I @VMODROOT/include
#include <dcimgui.h>
#include "backends/dcimgui_impl_glfw.h"
#include "backends/dcimgui_impl_vulkan.h"
pub const version = '1.91.9b'
pub const version_num = 19191
pub type C.ImFontBuilderIO = voidptr
pub type C.ImDrawListSharedData = voidptr
pub type C.ImGuiContext = voidptr
pub type C.va_list = voidptr
pub type C.ImGuiInputTextCallback = voidptr
pub type C.ImGuiSizeCallback = voidptr
pub type C.ImWchar = voidptr
pub type C.ImVec4 = voidptr

// THIS FILE HAS BEEN AUTO-GENERATED BY THE 'DEAR BINDINGS' GENERATOR.
// **DO NOT EDIT DIRECTLY**
// https://github.com/dearimgui/dear_bindings
// dear imgui, v1.91.9b
// (headers)
// Help:
// - See links below.
// - Call and read ImGui::ShowDemoWindow() in imgui_demo.cpp. All applications in examples/ are doing that.
// - Read top of imgui.cpp for more details, links and comments.
// - Add '#define IMGUI_DEFINE_MATH_OPERATORS' before including this file (or in imconfig.h) to access courtesy maths operators for ImVec2 and C.ImVec4.
// Resources:
// - FAQ ........................ https://dearimgui.com/faq (in repository as docs/FAQ.md)
// - Homepage ................... https://github.com/ocornut/imgui
// - Releases & changelog ....... https://github.com/ocornut/imgui/releases
// - Gallery .................... https://github.com/ocornut/imgui/issues?q=label%3Agallery (please post your screenshots/video there!)
// - Wiki ....................... https://github.com/ocornut/imgui/wiki (lots of good stuff there)
//   - Getting Started            https://github.com/ocornut/imgui/wiki/Getting-Started (how to integrate in an existing app by adding ~25 lines of code)
//   - Third-party Extensions     https://github.com/ocornut/imgui/wiki/Useful-Extensions (ImPlot & many more)
//   - Bindings/Backends          https://github.com/ocornut/imgui/wiki/Bindings (language bindings, backends for various tech/engines)
//   - Glossary                   https://github.com/ocornut/imgui/wiki/Glossary
//   - Debug Tools                https://github.com/ocornut/imgui/wiki/Debug-Tools
//   - Software using Dear ImGui  https://github.com/ocornut/imgui/wiki/Software-using-dear-imgui
// - Issues & support ........... https://github.com/ocornut/imgui/issues
// - Test Engine & Automation ... https://github.com/ocornut/imgui_test_engine (test suite, test engine to automate your apps)
// For first-time users having issues compiling/linking/running/loading fonts:
// please post in https://github.com/ocornut/imgui/discussions if you cannot find a solution in resources above.
// Everything else should be asked in 'Issues'! We are building a database of cross-linked knowledge there.
// Library Version
// (Integer encoded as XYYZZ for use in #if preprocessor conditionals, e.g. '#if IMGUI_VERSION_NUM >= 12345')
//
//
//Index of this file:
//// [SECTION] Header mess
//// [SECTION] Forward declarations and basic types
//// [SECTION] Texture identifier (ImTextureID)
//// [SECTION] Dear ImGui end-user API functions
//// [SECTION] Flags & Enumerations
//// [SECTION] Tables API flags and structures  TableFlags, TableColumnFlags, TableRowFlags, TableBgTarget, ImGuiTableSortSpecs, ImGuiTableColumnSortSpecs)
//// [SECTION] Helpers: Debug log, Memory allocations macros, ImVector<>
//// [SECTION] ImGuiStyle
//// [SECTION] ImGuiIO
//// [SECTION] Misc data structures (ImGuiInputTextCallbackData, ImGuiSizeCallbackData, ImGuiPayload)
//// [SECTION] Helpers  OnceUponAFrame, ImGuiTextFilter, ImGuiTextBuffer, ImGuiStorage, ImGuiListClipper, Math Operators, ImColor)
//// [SECTION] Multi-Select API flags and structures  MultiSelectFlags, ImGuiMultiSelectIO, ImGuiSelectionRequest, ImGuiSelectionBasicStorage, ImGuiSelectionExternalStorage)
//// [SECTION] Drawing API (ImDrawCallback, ImDrawCmd, ImDrawIdx, ImDrawVert, ImDrawChannel, ImDrawListSplitter, ImDrawFlags, ImDrawListFlags, ImDrawList, ImDrawData)
//// [SECTION] Font API (ImFontConfig, ImFontGlyph, ImFontGlyphRangesBuilder, ImFontAtlasFlags, ImFontAtlas, ImFont)
//// [SECTION] Viewports (ImGuiViewportFlags, ImGuiViewport)
//// [SECTION] ImGuiPlatformIO + other Platform Dependent Interfaces  PlatformImeData)
//// [SECTION] Obsolete functions and types
//
//
// Configuration file with compile-time options
// (edit imconfig.h or '#define IMGUI_USER_CONFIG "myfilename.h" from your build system)
// #ifdef IMGUI_USER_CONFIG
//-----------------------------------------------------------------------------
// [SECTION] Header mess
//-----------------------------------------------------------------------------
// Includes
// Define attributes of all API symbols declarations (e.g. for DLL under Windows)
// CIMGUI_API is used for core imgui functions, CIMGUI_IMPL_API is used for the default backends files (imgui_impl_xxx.h)
// Using dear imgui via a shared library is not recommended: we don't guarantee backward nor forward ABI compatibility + this is a call-heavy library and function call overhead adds up.
// #ifndef CIMGUI_API
// #ifndef CIMGUI_IMPL_API
// Helper Macros
// You can override the default assert handler by editing imconfig.h
// #ifndef IM_ASSERT
// Size of a static C-style array. Don't use on pointers!
// Used to silence "unused variable warnings". Often useful as asserts may be stripped out from final builds.
// Check that version and structures layouts are matching between compiled imgui code and caller. Read comments above DebugCheckVersionAndDataLayout() for details.
// Helper Macros - IM_FMTARGS, IM_FMTLIST: Apply printf-style warnings to our formatting functions.
// (MSVC provides an equivalent mechanism via SAL Annotations but it would require the macros in a different
//  location. e.g. #include <sal.h> + void myprintf(_Printf_format_string_ const char* format, ...))
// #if !defined(IMGUI_USE_STB_SPRINTF)&&(defined(__clang__)|| defined(__GNUC__))
// #if !defined(IMGUI_USE_STB_SPRINTF)&& defined(__MINGW32__)&&!defined(__clang__)
// Disable some of MSVC most aggressive Debug runtime checks in function header/footer (used in some simple/low-level functions)
// #if defined(_MSC_VER)&&!defined(__clang__)&&!defined(__INTEL_COMPILER)&&!defined(IMGUI_DEBUG_PARANOID)
// Warnings
// [Static Analyzer] Variable 'XXX' is uninitialized. Always initialize a member variable (type.6).
// #ifdef _MSC_VER
// warning: unknown warning group 'xxx'
// #if __has_warning("-Wunknown-warning-option")
// warning: unknown warning group 'xxx'
// warning: use of old-style cast
// warning: comparing floating point with == or != is unsafe
// warning: zero as null pointer constant
// warning: identifier '_Xxx' is reserved because it starts with '_' followed by a capital letter
// warning: 'xxx' is an unsafe pointer used for buffer access
// warning: first argument in call to 'memset' is a pointer to non-trivially copyable type
// warning: unknown option after '#pragma GCC diagnostic' kind
// warning: comparing floating-point with '==' or '!=' is unsafe
// [__GNUC__ >= 8] warning: 'memset/memcpy' clearing/writing an object of type 'xxxx' with no trivial copy-assignment; use assignment or value-initialization instead
// #if defined(__GNUC__)
// #if defined(__clang__)
//-----------------------------------------------------------------------------
// [SECTION] Forward declarations and basic types
// Auto-generated forward declarations for C header
// ImDrawIdx: vertex index. [Compile-time configurable type]
// - To use 16-bit indices + allow large meshes: backend need to set 'io.BackendFlags |= BackendFlags_RendererHasVtxOffset' and handle ImDrawCmd::VtxOffset (recommended).
// - To use 32-bit indices: override with '#define ImDrawIdx unsigned int' in your imconfig.h file.
type ImDrawIdx = u16
// Default: 16-bit (for maximum compatibility with renderer backends)
// #ifndef ImDrawIdx
//-----------------------------------------------------------------------------
// Scalar data types
type ID = u32
// A unique ID used by widgets (typically the result of hashing a stack of string)
type ImS8 = i8
// 8-bit signed integer
type ImU8 = u8
// 8-bit unsigned integer
type ImS16 = i16
// 16-bit signed integer
type ImU16 = u16
// 16-bit unsigned integer
type ImS32 = int
// 32-bit signed integer == int
type ImU32 = u32
// 32-bit unsigned integer (often used to store packed colors)
type ImS64 = i64
// 64-bit signed integer
type ImU64 = i64
// 64-bit unsigned integer
// Forward declarations: ImDrawList, ImFontAtlas layer
// Temporary storage to output draw commands out of order, used by ImDrawListSplitter and ImDrawList::ChannelsSplit()
// A single draw command within a parent ImDrawList (generally maps to 1 GPU draw call, unless it is a callback)
// All draw command lists required to render the frame + pos/size coordinates to use for the projection matrix.
// A single draw command list (generally one per window, conceptually you may see this as a dynamic "mesh" builder)
// Data shared among multiple draw lists (typically owned by parent ImGui context, but you may create one yourself)
// Helper to split a draw list into different layers which can be drawn into out of order, then flattened back.
// A single vertex (pos + uv + col = 20 bytes by default. Override layout with IMGUI_OVERRIDE_DRAWVERT_STRUCT_LAYOUT)
// Runtime data for a single font within a parent ImFontAtlas
// Runtime data for multiple fonts, bake multiple fonts into a single texture, TTF/OTF font loader
// Opaque interface to a font builder (stb_truetype or FreeType).
// Configuration data when adding a font or merging fonts
// A single font glyph (code point + coordinates within in ImFontAtlas + offset)
// Helper to build glyph ranges from text/string data
// Helper functions to create a color that can be converted to either u32 or float4 (*OBSOLETE* please avoid using)
// Forward declarations: ImGui layer
// Dear ImGui context (opaque structure, unless including imgui_internal.h)
// Main configuration and I/O between your application and ImGui (also see: ImGuiPlatformIO)
// Shared state of InputText() when using custom C.ImGuiInputTextCallback (rare/advanced use)
// Storage for ImGuiIO and IsKeyDown(), IsKeyPressed() etc functions.
// Helper to manually clip large list of items
// Structure to interact with a BeginMultiSelect()/EndMultiSelect() block
// User data payload for drag and drop operations
// Interface between platform/renderer backends and ImGui (e.g. Clipboard, IME hooks). Extends ImGuiIO. In docking branch, this gets extended to support multi-viewports.
// Platform IME data for io.PlatformSetImeDataFn() function.
// Optional helper to store multi-selection state + apply multi-selection requests.
//Optional helper to apply multi-selection requests to existing randomly accessible storage.
// A selection request (stored in ImGuiMultiSelectIO)
// Callback data when using SetNextWindowSizeConstraints() (rare/advanced use)
// Helper for key->value storage (container sorted by key)
// Helper for key->value storage (pair)
// Runtime data for styling/colors
// Sorting specifications for a table (often handling sort specs for a single column, occasionally more)
// Sorting specification for one column of a table
// Helper to hold and append into a text buffer (~string builder)
// Helper to parse and apply text filters (e.g. "aaaaa[,bbbbb][,ccccc]")
// A Platform Window (always only one in 'master' branch), in the future may represent Platform Monitor
// Enumerations
// - We don't use strongly typed enums much because they add constraints (can't extend in private code, can't store typed in bit fields, extra casting on iteration)
// - Tip: Use your programming IDE navigation facilities on the names in the _central column_ below to find the actual flags/enum lists!
//   - In Visual Studio: CTRL+comma ("Edit.GoToAll") can follow symbols inside comments, whereas CTRL+F12 ("Edit.GoToImplementation") cannot.
//   - In Visual Studio w/ Visual Assist installed: ALT+G ("VAssistX.GoToImplementation") can also follow symbols inside comments.
//   - In VS Code, CLion, etc.: CTRL+click can follow symbols inside comments.
type Dir = int
// -> enum Dir              // Enum: A cardinal direction (Left, Right, Up, Down)
type Key = int
// -> enum Key              // Enum: A key identifier  Key_XXX or Mod_XXX value)
type MouseSource = int
// -> enum MouseSource      // Enum; A mouse input source identifier (Mouse, TouchScreen, Pen)
type SortDirection = u8
// -> enum SortDirection    // Enum: A sorting direction (ascending or descending)
type Col = int
// -> enum Col_             // Enum: A color identifier for styling
type Cond = int
// -> enum Cond_            // Enum: A condition for many Set*() functions
type DataType = int
// -> enum DataType_        // Enum: A primary data type
type MouseButton = int
// -> enum MouseButton_     // Enum: A mouse button identifier (0=left, 1=right, 2=middle)
type MouseCursor = int
// -> enum MouseCursor_     // Enum: A mouse cursor shape
type ImGuiStyleVar = int
// -> enum ImGuiStyleVar_        // Enum: A variable identifier for styling
type TableBgTarget = int
// -> enum TableBgTarget_   // Enum: A color target for TableSetBgColor()
// Flags (declared as int to allow using as flags without overhead, and to not pollute the top of this file)
// - Tip: Use your programming IDE navigation facilities on the names in the _central column_ below to find the actual flags/enum lists!
//   - In Visual Studio: CTRL+comma ("Edit.GoToAll") can follow symbols inside comments, whereas CTRL+F12 ("Edit.GoToImplementation") cannot.
//   - In Visual Studio w/ Visual Assist installed: ALT+G ("VAssistX.GoToImplementation") can also follow symbols inside comments.
//   - In VS Code, CLion, etc.: CTRL+click can follow symbols inside comments.
type ImDrawFlags = int
// -> enum ImDrawFlags_          // Flags: for ImDrawList functions
type ImDrawListFlags = int
// -> enum ImDrawListFlags_      // Flags: for ImDrawList instance
type ImFontAtlasFlags = int
// -> enum ImFontAtlasFlags_     // Flags: for ImFontAtlas build
type BackendFlags = int
// -> enum BackendFlags_    // Flags: for io.BackendFlags
type ButtonFlags = int
// -> enum ButtonFlags_     // Flags: for InvisibleButton()
type ChildFlags = int
// -> enum ChildFlags_      // Flags: for BeginChild()
type ColorEditFlags = int
// -> enum ColorEditFlags_  // Flags: for ColorEdit4(), ColorPicker4() etc.
type ConfigFlags = int
// -> enum ConfigFlags_     // Flags: for io.ConfigFlags
type ComboFlags = int
// -> enum ComboFlags_      // Flags: for BeginCombo()
type DragDropFlags = int
// -> enum DragDropFlags_   // Flags: for BeginDragDropSource(), AcceptDragDropPayload()
type FocusedFlags = int
// -> enum FocusedFlags_    // Flags: for IsWindowFocused()
type HoveredFlags = int
// -> enum HoveredFlags_    // Flags: for IsItemHovered(), IsWindowHovered() etc.
type InputFlags = int
// -> enum InputFlags_      // Flags: for Shortcut(), SetNextItemShortcut()
type InputTextFlags = int
// -> enum InputTextFlags_  // Flags: for InputText(), InputTextMultiline()
type ItemFlags = int
// -> enum ItemFlags_       // Flags: for PushItemFlag(), shared by all items
type KeyChord = int
// -> Key | Mod_XXX    // Flags: for IsKeyChordPressed(), Shortcut() etc. an Key optionally OR-ed with one or more Mod_XXX values.
type PopupFlags = int
// -> enum PopupFlags_      // Flags: for OpenPopup*(), BeginPopupContext*(), IsPopupOpen()
type MultiSelectFlags = int
// -> enum MultiSelectFlags_// Flags: for BeginMultiSelect()
type SelectableFlags = int
// -> enum SelectableFlags_ // Flags: for Selectable()
type SliderFlags = int
// -> enum SliderFlags_     // Flags: for DragFloat(), DragInt(), SliderFloat(), SliderInt() etc.
type TabBarFlags = int
// -> enum TabBarFlags_     // Flags: for BeginTabBar()
type TabItemFlags = int
// -> enum TabItemFlags_    // Flags: for BeginTabItem()
type TableFlags = int
// -> enum TableFlags_      // Flags: For BeginTable()
type TableColumnFlags = int
// -> enum TableColumnFlags_// Flags: For TableSetupColumn()
type TableRowFlags = int
// -> enum TableRowFlags_   // Flags: For TableNextRow()
type TreeNodeFlags = int
// -> enum TreeNodeFlags_   // Flags: for TreeNode(), TreeNodeEx(), CollapsingHeader()
type ImGuiViewportFlags = int
// -> enum ImGuiViewportFlags_   // Flags: for ImGuiViewport
type WindowFlags = int
// -> enum WindowFlags_     // Flags: for Begin(), BeginChild()
// Character types
// (we generally use UTF-8 encoded string in the API. This is storage specifically for a decoded character used for keyboard input and display)
type ImWchar32 = u32
// A single decoded U32 character/code point. We encode them as multi bytes UTF-8 when used in strings.
type ImWchar16 = u16
// A single decoded U16 character/code point. We encode them as multi bytes UTF-8 when used in strings.
// C.ImWchar [configurable type: override in imconfig.h with '#define IMGUI_USE_WCHAR32' to support Unicode planes 1-16]
// Multi-Selection item index or identifier when using BeginMultiSelect()
// - Used by SetNextItemSelectionUserData() + and inside ImGuiMultiSelectIO structure.
// - Most users are likely to use this store an item INDEX but this may be used to store a POINTER/ID as well. Read comments near ImGuiMultiSelectIO for details.
type SelectionUserData = i64
// Callback and functions types
// Callback function for ImGui::InputText()
// Callback function for ImGui::SetNextWindowSizeConstraints()
type MemAllocFunc = fn (usize, voidptr) voidptr
// Function signature for ImGui::SetAllocatorFunctions()
type MemFreeFunc = fn (voidptr, voidptr)
// Function signature for ImGui::SetAllocatorFunctions()
// ImVec2: 2D vector used to store positions, sizes etc. [Compile-time configurable type]
// - This is a frequently used type in the API. Consider using IM_VEC2_CLASS_EXTRA to create implicit cast from/to our preferred type.
// - Add '#define IMGUI_DEFINE_MATH_OPERATORS' before including this file (or in imconfig.h) to access courtesy maths operators for ImVec2 and C.ImVec4.
struct ImVec2 { 
	x f32
	y f32
}
// C.ImVec4: 4D vector used to store clipping rectangles, colors etc. [Compile-time configurable type]
struct ImTextureID { 
	x f32
	y f32
	z f32
	w f32
}
//-----------------------------------------------------------------------------
// [SECTION] Texture identifier (ImTextureID)
//-----------------------------------------------------------------------------
// ImTexture: user data for renderer backend to identify a texture [Compile-time configurable type]
// - To use something else than an opaque void* pointer: override with e.g. '#define ImTextureID MyTextureType*' in your imconfig.h file.
// - This can be whatever to you want it to be! read the FAQ about ImTextureID for details.
// - You can make this a structure with various constructors if you need. You will have to implement ==/!= operators.
// - (note: before v1.91.4 (2024/10/08) the default type for ImTextureID was void*. Use intermediary intptr_t cast and read FAQ if you have casting warnings)
// Default: store a pointer or an integer fitting in a pointer (most renderer backends are ok with that)
// #ifndef ImTextureID
//-----------------------------------------------------------------------------
// [SECTION] Dear ImGui end-user API functions
// (Note that ImGui:: being a namespace, you can add extra ImGui:: functions in your own separate file. Please don't modify imgui source files!)
//-----------------------------------------------------------------------------
// Context creation and access
// - Each context create its own ImFontAtlas by default. You may instance one yourself and pass it to CreateContext() to share a font atlas between contexts.
// - DLL users: heaps and globals are not shared across DLL boundaries! You will need to call SetCurrentContext() + SetAllocatorFunctions()
//   for each static/DLL boundary you are calling from. Read "Context and Memory Allocators" section of imgui.cpp for details.
@[c:'ImGui_CreateContext']
fn create_context(shared_font_atlas &ImFontAtlas) &C.ImGuiContext

@[c:'ImGui_DestroyContext']
fn destroy_context(ctx &C.ImGuiContext)

// NULL = destroy current context
@[c:'ImGui_GetCurrentContext']
fn get_current_context() &C.ImGuiContext

@[c:'ImGui_SetCurrentContext']
fn set_current_context(ctx &C.ImGuiContext)

// Main
@[c:'ImGui_GetIO']
fn get_io() &ImGuiIO

// access the ImGuiIO structure (mouse/keyboard/gamepad inputs, time, various configuration options/flags)
@[c:'ImGui_GetPlatformIO']
fn get_platform_io() &ImGuiPlatformIO

// access the ImGuiPlatformIO structure (mostly hooks/functions to connect to platform/renderer and OS Clipboard, IME etc.)
@[c:'ImGui_GetStyle']
fn get_style() &ImGuiStyle

// access the Style structure (colors, sizes). Always use PushStyleColor(), PushStyleVar() to modify style mid-frame!
@[c:'ImGui_NewFrame']
fn new_frame()

// start a new Dear ImGui frame, you can submit any command from this point until Render()/EndFrame().
@[c:'ImGui_EndFrame']
fn end_frame()

// ends the Dear ImGui frame. automatically called by Render(). If you don't need to render data (skipping rendering) you may call EndFrame() without Render()... but you'll have wasted CPU already! If you don't need to render, better to not create any windows and not call NewFrame() at all!
@[c:'ImGui_Render']
fn render()

// ends the Dear ImGui frame, finalize the draw data. You can then get call GetDrawData().
@[c:'ImGui_GetDrawData']
fn get_draw_data() &ImDrawData

// valid after Render() and until the next call to NewFrame(). this is what you have to render.
// Demo, Debug, Information
@[c:'ImGui_ShowDemoWindow']
fn show_demo_window(p_open &bool)

// create Demo window. demonstrate most ImGui features. call this to learn about the library! try to make it always available in your application!
@[c:'ImGui_ShowMetricsWindow']
fn show_metrics_window(p_open &bool)

// create Metrics/Debugger window. display Dear ImGui internals: windows, draw commands, various internal state, etc.
@[c:'ImGui_ShowDebugLogWindow']
fn show_debug_log_window(p_open &bool)

// create Debug Log window. display a simplified log of important dear imgui events.
@[c:'ImGui_ShowIDStackToolWindow']
fn show_ids_tack_tool_window()

// Implied p_open = NULL
@[c:'ImGui_ShowIDStackToolWindowEx']
fn show_ids_tack_tool_window_ex(p_open &bool)

// create Stack Tool window. hover items with mouse to query information about the source of their unique ID.
@[c:'ImGui_ShowAboutWindow']
fn show_about_window(p_open &bool)

// create About window. display Dear ImGui version, credits and build/system information.
@[c:'ImGui_ShowStyleEditor']
fn show_style_editor(ref &ImGuiStyle)

// add style editor block (not a window). you can pass in a reference ImGuiStyle structure to compare to, revert to and save to (else it uses the default style)
@[c:'ImGui_ShowStyleSelector']
fn show_style_selector(label &i8) bool

// add style selector block (not a window), essentially a combo listing the default styles.
@[c:'ImGui_ShowFontSelector']
fn show_font_selector(label &i8)

// add font selector block (not a window), essentially a combo listing the loaded fonts.
@[c:'ImGui_ShowUserGuide']
fn show_user_guide()

// add basic help/info block (not a window): how to manipulate ImGui as an end-user (mouse/keyboard controls).
@[c:'ImGui_GetVersion']
fn get_version() &i8

// get the compiled version string e.g. "1.80 WIP" (essentially the value for IMGUI_VERSION from the compiled version of imgui.cpp)
// Styles
@[c:'ImGui_StyleColorsDark']
fn style_colors_dark(dst &ImGuiStyle)

// new, recommended style (default)
@[c:'ImGui_StyleColorsLight']
fn style_colors_light(dst &ImGuiStyle)

// best used with borders and a custom, thicker font
@[c:'ImGui_StyleColorsClassic']
fn style_colors_classic(dst &ImGuiStyle)

// classic imgui style
// Windows
// - Begin() = push window to the stack and start appending to it. End() = pop window from the stack.
// - Passing 'bool* p_open != NULL' shows a window-closing widget in the upper-right corner of the window,
//   which clicking will set the boolean to false when clicked.
// - You may append multiple times to the same window during the same frame by calling Begin()/End() pairs multiple times.
//   Some information such as 'flags' or 'p_open' will only be considered by the first call to Begin().
// - Begin() return false to indicate the window is collapsed or fully clipped, so you may early out and omit submitting
//   anything to the window. Always call a matching End() for each Begin() call, regardless of its return value!
//   [Important: due to legacy reason, Begin/End and BeginChild/EndChild are inconsistent with all other functions
//    such as BeginMenu/EndMenu, BeginPopup/EndPopup, etc. where the EndXXX call should only be called if the corresponding
//    BeginXXX function returned true. Begin and BeginChild are the only odd ones out. Will be fixed in a future update.]
// - Note that the bottom of window stack always contains a window called "Debug".
@[c:'ImGui_Begin']
fn begin(name &i8, p_open &bool, flags WindowFlags) bool

@[c:'ImGui_End']
fn end()

// Child Windows
// - Use child windows to begin into a self-contained independent scrolling/clipping regions within a host window. Child windows can embed their own child.
// - Before 1.90 (November 2023), the  ChildFlags child_flags = 0" parameter was "bool border = false".
//   This API is backward compatible with old code, as we guarantee that ChildFlags_Borders == true.
//   Consider updating your old code:
//      BeginChild("Name", size, false)   -> Begin("Name", size, 0); or Begin("Name", size, ChildFlags_None);
//      BeginChild("Name", size, true)    -> Begin("Name", size, ChildFlags_Borders);
// - Manual sizing (each axis can use a different setting e.g. ImVec2(0.0f, 400.0f)):
//     == 0.0f: use remaining parent window size for this axis.
//      > 0.0f: use specified size for this axis.
//      < 0.0f: right/bottom-align to specified distance from available content boundaries.
// - Specifying ChildFlags_AutoResizeX or ChildFlags_AutoResizeY makes the sizing automatic based on child contents.
//   Combining both ChildFlags_AutoResizeX _and_ ChildFlags_AutoResizeY defeats purpose of a scrolling region and is NOT recommended.
// - BeginChild() returns false to indicate the window is collapsed or fully clipped, so you may early out and omit submitting
//   anything to the window. Always call a matching EndChild() for each BeginChild() call, regardless of its return value.
//   [Important: due to legacy reason, Begin/End and BeginChild/EndChild are inconsistent with all other functions
//    such as BeginMenu/EndMenu, BeginPopup/EndPopup, etc. where the EndXXX call should only be called if the corresponding
//    BeginXXX function returned true. Begin and BeginChild are the only odd ones out. Will be fixed in a future update.]
@[c:'ImGui_BeginChild']
fn begin_child(str_id &i8, size ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c:'ImGui_BeginChildID']
fn begin_child_id(id ID, size ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c:'ImGui_EndChild']
fn end_child()

// Windows Utilities
// - 'current window' = the window we are appending into while inside a Begin()/End() block. 'next window' = next window we will Begin() into.
@[c:'ImGui_IsWindowAppearing']
fn is_window_appearing() bool

@[c:'ImGui_IsWindowCollapsed']
fn is_window_collapsed() bool

@[c:'ImGui_IsWindowFocused']
fn is_window_focused(flags FocusedFlags) bool

// is current window focused? or its root/child, depending on flags. see flags for options.
@[c:'ImGui_IsWindowHovered']
fn is_window_hovered(flags HoveredFlags) bool

// is current window hovered and hoverable (e.g. not blocked by a popup/modal)? See HoveredFlags_ for options. IMPORTANT: If you are trying to check whether your mouse should be dispatched to Dear ImGui or to your underlying app, you should not use this function! Use the 'io.WantCaptureMouse' boolean for that! Refer to FAQ entry "How can I tell whether to dispatch mouse/keyboard to Dear ImGui or my application?" for details.
@[c:'ImGui_GetWindowDrawList']
fn get_window_draw_list() &ImDrawList

// get draw list associated to the current window, to append your own drawing primitives
@[c:'ImGui_GetWindowPos']
fn get_window_pos() ImVec2

// get current window position in screen space (IT IS UNLIKELY YOU EVER NEED TO USE THIS. Consider always using GetCursorScreenPos() and GetContentRegionAvail() instead)
@[c:'ImGui_GetWindowSize']
fn get_window_size() ImVec2

// get current window size (IT IS UNLIKELY YOU EVER NEED TO USE THIS. Consider always using GetCursorScreenPos() and GetContentRegionAvail() instead)
@[c:'ImGui_GetWindowWidth']
fn get_window_width() f32

// get current window width (IT IS UNLIKELY YOU EVER NEED TO USE THIS). Shortcut for GetWindowSize().x.
@[c:'ImGui_GetWindowHeight']
fn get_window_height() f32

// get current window height (IT IS UNLIKELY YOU EVER NEED TO USE THIS). Shortcut for GetWindowSize().y.
// Window manipulation
// - Prefer using SetNextXXX functions (before Begin) rather that SetXXX functions (after Begin).
@[c:'ImGui_SetNextWindowPos']
fn set_next_window_pos(pos ImVec2, cond Cond)

// Implied pivot = ImVec2(0, 0)
@[c:'ImGui_SetNextWindowPosEx']
fn set_next_window_pos_ex(pos ImVec2, cond Cond, pivot ImVec2)

// set next window position. call before Begin(). use pivot=(0.5f,0.5f) to center on given point, etc.
@[c:'ImGui_SetNextWindowSize']
fn set_next_window_size(size ImVec2, cond Cond)

// set next window size. set axis to 0.0f to force an auto-fit on this axis. call before Begin()
@[c:'ImGui_SetNextWindowSizeConstraints']
fn set_next_window_size_constraints(size_min ImVec2, size_max ImVec2, custom_callback C.ImGuiSizeCallback, custom_callback_data voidptr)

// set next window size limits. use 0.0f or FLT_MAX if you don't want limits. Use -1 for both min and max of same axis to preserve current size (which itself is a constraint). Use callback to apply non-trivial programmatic constraints.
@[c:'ImGui_SetNextWindowContentSize']
fn set_next_window_content_size(size ImVec2)

// set next window content size (~ scrollable client area, which enforce the range of scrollbars). Not including window decorations (title bar, menu bar, etc.) nor WindowPadding. set an axis to 0.0f to leave it automatic. call before Begin()
@[c:'ImGui_SetNextWindowCollapsed']
fn set_next_window_collapsed(collapsed bool, cond Cond)

// set next window collapsed state. call before Begin()
@[c:'ImGui_SetNextWindowFocus']
fn set_next_window_focus()

// set next window to be focused / top-most. call before Begin()
@[c:'ImGui_SetNextWindowScroll']
fn set_next_window_scroll(scroll ImVec2)

// set next window scrolling value (use < 0.0f to not affect a given axis).
@[c:'ImGui_SetNextWindowBgAlpha']
fn set_next_window_bg_alpha(alpha f32)

// set next window background color alpha. helper to easily override the Alpha component of Col_WindowBg/ChildBg/PopupBg. you may also use WindowFlags_NoBackground.
@[c:'ImGui_SetWindowPos']
fn set_window_pos(pos ImVec2, cond Cond)

// (not recommended) set current window position - call within Begin()/End(). prefer using SetNextWindowPos(), as this may incur tearing and side-effects.
@[c:'ImGui_SetWindowSize']
fn set_window_size(size ImVec2, cond Cond)

// (not recommended) set current window size - call within Begin()/End(). set to ImVec2(0, 0) to force an auto-fit. prefer using SetNextWindowSize(), as this may incur tearing and minor side-effects.
@[c:'ImGui_SetWindowCollapsed']
fn set_window_collapsed(collapsed bool, cond Cond)

// (not recommended) set current window collapsed state. prefer using SetNextWindowCollapsed().
@[c:'ImGui_SetWindowFocus']
fn set_window_focus()

// (not recommended) set current window to be focused / top-most. prefer using SetNextWindowFocus().
@[c:'ImGui_SetWindowFontScale']
fn set_window_font_scale(scale f32)

// [OBSOLETE] set font scale. Adjust IO.FontGlobalScale if you want to scale all windows. This is an old API! For correct scaling, prefer to reload font + rebuild ImFontAtlas + call style.ScaleAllSizes().
@[c:'ImGui_SetWindowPosStr']
fn set_window_pos_str(name &i8, pos ImVec2, cond Cond)

// set named window position.
@[c:'ImGui_SetWindowSizeStr']
fn set_window_size_str(name &i8, size ImVec2, cond Cond)

// set named window size. set axis to 0.0f to force an auto-fit on this axis.
@[c:'ImGui_SetWindowCollapsedStr']
fn set_window_collapsed_str(name &i8, collapsed bool, cond Cond)

// set named window collapsed state
@[c:'ImGui_SetWindowFocusStr']
fn set_window_focus_str(name &i8)

// set named window to be focused / top-most. use NULL to remove focus.
// Windows Scrolling
// - Any change of Scroll will be applied at the beginning of next frame in the first call to Begin().
// - You may instead use SetNextWindowScroll() prior to calling Begin() to avoid this delay, as an alternative to using SetScrollX()/SetScrollY().
@[c:'ImGui_GetScrollX']
fn get_scroll_x() f32

// get scrolling amount [0 .. GetScrollMaxX()]
@[c:'ImGui_GetScrollY']
fn get_scroll_y() f32

// get scrolling amount [0 .. GetScrollMaxY()]
@[c:'ImGui_SetScrollX']
fn set_scroll_x(scroll_x f32)

// set scrolling amount [0 .. GetScrollMaxX()]
@[c:'ImGui_SetScrollY']
fn set_scroll_y(scroll_y f32)

// set scrolling amount [0 .. GetScrollMaxY()]
@[c:'ImGui_GetScrollMaxX']
fn get_scroll_max_x() f32

// get maximum scrolling amount ~~ ContentSize.x - WindowSize.x - DecorationsSize.x
@[c:'ImGui_GetScrollMaxY']
fn get_scroll_max_y() f32

// get maximum scrolling amount ~~ ContentSize.y - WindowSize.y - DecorationsSize.y
@[c:'ImGui_SetScrollHereX']
fn set_scroll_here_x(center_x_ratio f32)

// adjust scrolling amount to make current cursor position visible. center_x_ratio=0.0: left, 0.5: center, 1.0: right. When using to make a "default/current item" visible, consider using SetItemDefaultFocus() instead.
@[c:'ImGui_SetScrollHereY']
fn set_scroll_here_y(center_y_ratio f32)

// adjust scrolling amount to make current cursor position visible. center_y_ratio=0.0: top, 0.5: center, 1.0: bottom. When using to make a "default/current item" visible, consider using SetItemDefaultFocus() instead.
@[c:'ImGui_SetScrollFromPosX']
fn set_scroll_from_pos_x(local_x f32, center_x_ratio f32)

// adjust scrolling amount to make given position visible. Generally GetCursorStartPos() + offset to compute a valid position.
@[c:'ImGui_SetScrollFromPosY']
fn set_scroll_from_pos_y(local_y f32, center_y_ratio f32)

// adjust scrolling amount to make given position visible. Generally GetCursorStartPos() + offset to compute a valid position.
// Parameters stacks (shared)
@[c:'ImGui_PushFont']
fn push_font(font &ImFont)

// use NULL as a shortcut to push default font
@[c:'ImGui_PopFont']
fn pop_font()

@[c:'ImGui_PushStyleColor']
fn push_style_color(idx Col, col ImU32)

// modify a style color. always use this if you modify the style after NewFrame().
@[c:'ImGui_PushStyleColorImVec4']
fn push_style_color_im_vec4(idx Col, col C.ImVec4)

@[c:'ImGui_PopStyleColor']
fn pop_style_color()

// Implied count = 1
@[c:'ImGui_PopStyleColorEx']
fn pop_style_color_ex(count int)

@[c:'ImGui_PushStyleVar']
fn push_style_var(idx ImGuiStyleVar, val f32)

// modify a style float variable. always use this if you modify the style after NewFrame()!
@[c:'ImGui_PushStyleVarImVec2']
fn push_style_var_im_vec2(idx ImGuiStyleVar, val ImVec2)

// modify a style ImVec2 variable. "
@[c:'ImGui_PushStyleVarX']
fn push_style_var_x(idx ImGuiStyleVar, val_x f32)

// modify X component of a style ImVec2 variable. "
@[c:'ImGui_PushStyleVarY']
fn push_style_var_y(idx ImGuiStyleVar, val_y f32)

// modify Y component of a style ImVec2 variable. "
@[c:'ImGui_PopStyleVar']
fn pop_style_var()

// Implied count = 1
@[c:'ImGui_PopStyleVarEx']
fn pop_style_var_ex(count int)

@[c:'ImGui_PushItemFlag']
fn push_item_flag(option ItemFlags, enabled bool)

// modify specified shared item flag, e.g. PushItemFlag ItemFlags_NoTabStop, true)
@[c:'ImGui_PopItemFlag']
fn pop_item_flag()

// Parameters stacks (current window)
@[c:'ImGui_PushItemWidth']
fn push_item_width(item_width f32)

// push width of items for common large "item+label" widgets. >0.0f: width in pixels, <0.0f align xx pixels to the right of window (so -FLT_MIN always align width to the right side).
@[c:'ImGui_PopItemWidth']
fn pop_item_width()

@[c:'ImGui_SetNextItemWidth']
fn set_next_item_width(item_width f32)

// set width of the _next_ common large "item+label" widget. >0.0f: width in pixels, <0.0f align xx pixels to the right of window (so -FLT_MIN always align width to the right side)
@[c:'ImGui_CalcItemWidth']
fn calc_item_width() f32

// width of item given pushed settings and current cursor position. NOT necessarily the width of last item unlike most 'Item' functions.
@[c:'ImGui_PushTextWrapPos']
fn push_text_wrap_pos(wrap_local_pos_x f32)

// push word-wrapping position for Text*() commands. < 0.0f: no wrapping; 0.0f: wrap to end of window (or column); > 0.0f: wrap at 'wrap_pos_x' position in window local space
@[c:'ImGui_PopTextWrapPos']
fn pop_text_wrap_pos()

// Style read access
// - Use the ShowStyleEditor() function to interactively see/edit the colors.
@[c:'ImGui_GetFont']
fn get_font() &ImFont

// get current font
@[c:'ImGui_GetFontSize']
fn get_font_size() f32

// get current font size (= height in pixels) of current font with current scale applied
@[c:'ImGui_GetFontTexUvWhitePixel']
fn get_font_tex_uv_white_pixel() ImVec2

// get UV coordinate for a white pixel, useful to draw custom shapes via the ImDrawList API
@[c:'ImGui_GetColorU32']
fn get_color_u32(idx Col) ImU32

// Implied alpha_mul = 1.0f
@[c:'ImGui_GetColorU32Ex']
fn get_color_u32_ex(idx Col, alpha_mul f32) ImU32

// retrieve given style color with style alpha applied and optional extra alpha multiplier, packed as a 32-bit value suitable for ImDrawList
@[c:'ImGui_GetColorU32ImVec4']
fn get_color_u32_im_vec4(col C.ImVec4) ImU32

// retrieve given color with style alpha applied, packed as a 32-bit value suitable for ImDrawList
@[c:'ImGui_GetColorU32ImU32']
fn get_color_u32_im_u32(col ImU32) ImU32

// Implied alpha_mul = 1.0f
@[c:'ImGui_GetColorU32ImU32Ex']
fn get_color_u32_im_u32_ex(col ImU32, alpha_mul f32) ImU32

// retrieve given color with style alpha applied, packed as a 32-bit value suitable for ImDrawList
@[c:'ImGui_GetStyleColorVec4']
fn get_style_color_vec4(idx Col) &C.ImVec4

// retrieve style color as stored in ImGuiStyle structure. use to feed back into PushStyleColor(), otherwise use GetColorU32() to get style color with style alpha baked in.
// Layout cursor positioning
// - By "cursor" we mean the current output position.
// - The typical widget behavior is to output themselves at the current cursor position, then move the cursor one line down.
// - You can call SameLine() between widgets to undo the last carriage return and output at the right of the preceding widget.
// - YOU CAN DO 99% OF WHAT YOU NEED WITH ONLY GetCursorScreenPos() and GetContentRegionAvail().
// - Attention! We currently have inconsistencies between window-local and absolute positions we will aim to fix with future API:
//    - Absolute coordinate:        GetCursorScreenPos(), SetCursorScreenPos(), all ImDrawList:: functions. -> this is the preferred way forward.
//    - Window-local coordinates:   SameLine(offset), GetCursorPos(), SetCursorPos(), GetCursorStartPos(), PushTextWrapPos()
//    - Window-local coordinates:   GetContentRegionMax(), GetWindowContentRegionMin(), GetWindowContentRegionMax() --> all obsoleted. YOU DON'T NEED THEM.
// - GetCursorScreenPos() = GetCursorPos() + GetWindowPos(). GetWindowPos() is almost only ever useful to convert from window-local to absolute coordinates. Try not to use it.
@[c:'ImGui_GetCursorScreenPos']
fn get_cursor_screen_pos() ImVec2

// cursor position, absolute coordinates. THIS IS YOUR BEST FRIEND (prefer using this rather than GetCursorPos(), also more useful to work with ImDrawList API).
@[c:'ImGui_SetCursorScreenPos']
fn set_cursor_screen_pos(pos ImVec2)

// cursor position, absolute coordinates. THIS IS YOUR BEST FRIEND.
@[c:'ImGui_GetContentRegionAvail']
fn get_content_region_avail() ImVec2

// available space from current position. THIS IS YOUR BEST FRIEND.
@[c:'ImGui_GetCursorPos']
fn get_cursor_pos() ImVec2

// [window-local] cursor position in window-local coordinates. This is not your best friend.
@[c:'ImGui_GetCursorPosX']
fn get_cursor_pos_x() f32

// [window-local] "
@[c:'ImGui_GetCursorPosY']
fn get_cursor_pos_y() f32

// [window-local] "
@[c:'ImGui_SetCursorPos']
fn set_cursor_pos(local_pos ImVec2)

// [window-local] "
@[c:'ImGui_SetCursorPosX']
fn set_cursor_pos_x(local_x f32)

// [window-local] "
@[c:'ImGui_SetCursorPosY']
fn set_cursor_pos_y(local_y f32)

// [window-local] "
@[c:'ImGui_GetCursorStartPos']
fn get_cursor_start_pos() ImVec2

// [window-local] initial cursor position, in window-local coordinates. Call GetCursorScreenPos() after Begin() to get the absolute coordinates version.
// Other layout functions
@[c:'ImGui_Separator']
fn separator()

// separator, generally horizontal. inside a menu bar or in horizontal layout mode, this becomes a vertical separator.
@[c:'ImGui_SameLine']
fn same_line()

// Implied offset_from_start_x = 0.0f, spacing = -1.0f
@[c:'ImGui_SameLineEx']
fn same_line_ex(offset_from_start_x f32, spacing f32)

// call between widgets or groups to layout them horizontally. X position given in window coordinates.
@[c:'ImGui_NewLine']
fn new_line()

// undo a SameLine() or force a new line when in a horizontal-layout context.
@[c:'ImGui_Spacing']
fn spacing()

// add vertical spacing.
@[c:'ImGui_Dummy']
fn dummy(size ImVec2)

// add a dummy item of given size. unlike InvisibleButton(), Dummy() won't take the mouse click or be navigable into.
@[c:'ImGui_Indent']
fn indent()

// Implied indent_w = 0.0f
@[c:'ImGui_IndentEx']
fn indent_ex(indent_w f32)

// move content position toward the right, by indent_w, or style.IndentSpacing if indent_w <= 0
@[c:'ImGui_Unindent']
fn unindent()

// Implied indent_w = 0.0f
@[c:'ImGui_UnindentEx']
fn unindent_ex(indent_w f32)

// move content position back to the left, by indent_w, or style.IndentSpacing if indent_w <= 0
@[c:'ImGui_BeginGroup']
fn begin_group()

// lock horizontal starting position
@[c:'ImGui_EndGroup']
fn end_group()

// unlock horizontal starting position + capture the whole group bounding box into one "item" (so you can use IsItemHovered() or layout primitives such as SameLine() on whole group, etc.)
@[c:'ImGui_AlignTextToFramePadding']
fn align_text_to_frame_padding()

// vertically align upcoming text baseline to FramePadding.y so that it will align properly to regularly framed items (call if you have text on a line before a framed item)
@[c:'ImGui_GetTextLineHeight']
fn get_text_line_height() f32

// ~ FontSize
@[c:'ImGui_GetTextLineHeightWithSpacing']
fn get_text_line_height_with_spacing() f32

// ~ FontSize + style.ItemSpacing.y (distance in pixels between 2 consecutive lines of text)
@[c:'ImGui_GetFrameHeight']
fn get_frame_height() f32

// ~ FontSize + style.FramePadding.y * 2
@[c:'ImGui_GetFrameHeightWithSpacing']
fn get_frame_height_with_spacing() f32

// ~ FontSize + style.FramePadding.y * 2 + style.ItemSpacing.y (distance in pixels between 2 consecutive lines of framed widgets)
// ID stack/scopes
// Read the FAQ (docs/FAQ.md or http://dearimgui.com/faq) for more details about how ID are handled in dear imgui.
// - Those questions are answered and impacted by understanding of the ID stack system:
//   - "Q: Why is my widget not reacting when I click on it?"
//   - "Q: How can I have widgets with an empty label?"
//   - "Q: How can I have multiple widgets with the same label?"
// - Short version: ID are hashes of the entire ID stack. If you are creating widgets in a loop you most likely
//   want to push a unique identifier (e.g. object pointer, loop index) to uniquely differentiate them.
// - You can also use the "Label##foobar" syntax within widget label to distinguish them from each others.
// - In this header file we use the "label"/"name" terminology to denote a string that will be displayed + used as an ID,
//   whereas "str_id" denote a string that is only used as an ID and not normally displayed.
@[c:'ImGui_PushID']
fn push_id(str_id &i8)

// push string into the ID stack (will hash string).
@[c:'ImGui_PushIDStr']
fn push_ids_tr(str_id_begin &i8, str_id_end &i8)

// push string into the ID stack (will hash string).
@[c:'ImGui_PushIDPtr']
fn push_idp_tr(ptr_id voidptr)

// push pointer into the ID stack (will hash pointer).
@[c:'ImGui_PushIDInt']
fn push_idi_nt(int_id int)

// push integer into the ID stack (will hash integer).
@[c:'ImGui_PopID']
fn pop_id()

// pop from the ID stack.
@[c:'ImGui_GetID']
fn get_id(str_id &i8) ID

// calculate unique ID (hash of whole ID stack + given parameter). e.g. if you want to query into ImGuiStorage yourself
@[c:'ImGui_GetIDStr']
fn get_ids_tr(str_id_begin &i8, str_id_end &i8) ID

@[c:'ImGui_GetIDPtr']
fn get_idp_tr(ptr_id voidptr) ID

@[c:'ImGui_GetIDInt']
fn get_idi_nt(int_id int) ID

// Widgets: Text
@[c:'ImGui_TextUnformatted']
fn text_unformatted(text &i8)

// Implied text_end = NULL
@[c:'ImGui_TextUnformattedEx']
fn text_unformatted_ex(text &i8, text_end &i8)

// raw text without formatting. Roughly equivalent to Text("%s", text) but: A) doesn't require null terminated string if 'text_end' is specified, B) it's faster, no memory copy is done, no buffer size limits, recommended for long chunks of text.
@[c2v_variadic]
@[c:'ImGui_Text']
fn text(fmt &i8)

// formatted text
@[c:'ImGui_TextV']
fn text_v(fmt &i8, args C.va_list)

@[c2v_variadic]
@[c:'ImGui_TextColored']
fn text_colored(col C.ImVec4, fmt &i8)

// shortcut for PushStyleColor Col_Text, col); Text(fmt, ...); PopStyleColor();
@[c:'ImGui_TextColoredV']
fn text_colored_v(col C.ImVec4, fmt &i8, args C.va_list)

@[c2v_variadic]
@[c:'ImGui_TextDisabled']
fn text_disabled(fmt &i8)

// shortcut for PushStyleColor Col_Text, style.Colors Col_TextDisabled]); Text(fmt, ...); PopStyleColor();
@[c:'ImGui_TextDisabledV']
fn text_disabled_v(fmt &i8, args C.va_list)

@[c2v_variadic]
@[c:'ImGui_TextWrapped']
fn text_wrapped(fmt &i8)

// shortcut for PushTextWrapPos(0.0f); Text(fmt, ...); PopTextWrapPos();. Note that this won't work on an auto-resizing window if there's no other widgets to extend the window width, yoy may need to set a size using SetNextWindowSize().
@[c:'ImGui_TextWrappedV']
fn text_wrapped_v(fmt &i8, args C.va_list)

@[c2v_variadic]
@[c:'ImGui_LabelText']
fn label_text(label &i8, fmt &i8)

// display text+label aligned the same way as value+label widgets
@[c:'ImGui_LabelTextV']
fn label_text_v(label &i8, fmt &i8, args C.va_list)

@[c2v_variadic]
@[c:'ImGui_BulletText']
fn bullet_text(fmt &i8)

// shortcut for Bullet()+Text()
@[c:'ImGui_BulletTextV']
fn bullet_text_v(fmt &i8, args C.va_list)

@[c:'ImGui_SeparatorText']
fn separator_text(label &i8)

// currently: formatted text with a horizontal line
// Widgets: Main
// - Most widgets return true when the value has been changed or when pressed/selected
// - You may also use one of the many IsItemXXX functions (e.g. IsItemActive, IsItemHovered, etc.) to query widget state.
@[c:'ImGui_Button']
fn button(label &i8) bool

// Implied size = ImVec2(0, 0)
@[c:'ImGui_ButtonEx']
fn button_ex(label &i8, size ImVec2) bool

// button
@[c:'ImGui_SmallButton']
fn small_button(label &i8) bool

// button with (FramePadding.y == 0) to easily embed within text
@[c:'ImGui_InvisibleButton']
fn invisible_button(str_id &i8, size ImVec2, flags ButtonFlags) bool

// flexible button behavior without the visuals, frequently useful to build custom behaviors using the public api (along with IsItemActive, IsItemHovered, etc.)
@[c:'ImGui_ArrowButton']
fn arrow_button(str_id &i8, dir Dir) bool

// square button with an arrow shape
@[c:'ImGui_Checkbox']
fn checkbox(label &i8, v &bool) bool

@[c:'ImGui_CheckboxFlagsIntPtr']
fn checkbox_flags_int_ptr(label &i8, flags &int, flags_value int) bool

@[c:'ImGui_CheckboxFlagsUintPtr']
fn checkbox_flags_uint_ptr(label &i8, flags &u32, flags_value u32) bool

@[c:'ImGui_RadioButton']
fn radio_button(label &i8, active bool) bool

// use with e.g. if (RadioButton("one", my_value==1)) { my_value = 1; }
@[c:'ImGui_RadioButtonIntPtr']
fn radio_button_int_ptr(label &i8, v &int, v_button int) bool

// shortcut to handle the above pattern when value is an integer
@[c:'ImGui_ProgressBar']
fn progress_bar(fraction f32, size_arg ImVec2, overlay &i8)

@[c:'ImGui_Bullet']
fn bullet()

// draw a small circle + keep the cursor on the same line. advance cursor x position by GetTreeNodeToLabelSpacing(), same distance that TreeNode() uses
@[c:'ImGui_TextLink']
fn text_link(label &i8) bool

// hyperlink text button, return true when clicked
@[c:'ImGui_TextLinkOpenURL']
fn text_link_open_url(label &i8)

// Implied url = NULL
@[c:'ImGui_TextLinkOpenURLEx']
fn text_link_open_urle_x(label &i8, url &i8)

// hyperlink text button, automatically open file/url when clicked
// Widgets: Images
// - Read about ImTextureID here: https://github.com/ocornut/imgui/wiki/Image-Loading-and-Displaying-Examples
// - 'uv0' and 'uv1' are texture coordinates. Read about them from the same link above.
// - Image() pads adds style.ImageBorderSize on each side, ImageButton() adds style.FramePadding on each side.
// - ImageButton() draws a background based on regular Button() color + optionally an inner background if specified.
@[c:'ImGui_Image']
fn image(user_texture_id ImTextureID, image_size ImVec2)

// Implied uv0 = ImVec2(0, 0), uv1 = ImVec2(1, 1)
@[c:'ImGui_ImageEx']
fn image_ex(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2)

@[c:'ImGui_ImageWithBg']
fn image_with_bg(user_texture_id ImTextureID, image_size ImVec2)

// Implied uv0 = ImVec2(0, 0), uv1 = ImVec2(1, 1), bg_col = C.ImVec4(0, 0, 0, 0), tint_col = C.ImVec4(1, 1, 1, 1)
@[c:'ImGui_ImageWithBgEx']
fn image_with_bg_ex(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col C.ImVec4, tint_col C.ImVec4)

@[c:'ImGui_ImageButton']
fn image_button(str_id &i8, user_texture_id ImTextureID, image_size ImVec2) bool

// Implied uv0 = ImVec2(0, 0), uv1 = ImVec2(1, 1), bg_col = C.ImVec4(0, 0, 0, 0), tint_col = C.ImVec4(1, 1, 1, 1)
@[c:'ImGui_ImageButtonEx']
fn image_button_ex(str_id &i8, user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col C.ImVec4, tint_col C.ImVec4) bool

// Widgets: Combo Box (Dropdown)
// - The BeginCombo()/EndCombo() api allows you to manage your contents and selection state however you want it, by creating e.g. Selectable() items.
// - The old Combo() api are helpers over BeginCombo()/EndCombo() which are kept available for convenience purpose. This is analogous to how ListBox are created.
@[c:'ImGui_BeginCombo']
fn begin_combo(label &i8, preview_value &i8, flags ComboFlags) bool

@[c:'ImGui_EndCombo']
fn end_combo()

// only call EndCombo() if BeginCombo() returns true!
@[c:'ImGui_ComboChar']
fn combo_char(label &i8, current_item &int, items &&u8, items_count int) bool

// Implied popup_max_height_in_items = -1
@[c:'ImGui_ComboCharEx']
fn combo_char_ex(label &i8, current_item &int, items &&u8, items_count int, popup_max_height_in_items int) bool

@[c:'ImGui_Combo']
fn combo(label &i8, current_item &int, items_separated_by_zeros &i8) bool

// Implied popup_max_height_in_items = -1
@[c:'ImGui_ComboEx']
fn combo_ex(label &i8, current_item &int, items_separated_by_zeros &i8, popup_max_height_in_items int) bool

// Separate items with \0 within a string, end item-list with \0\0. e.g. "One\0Two\0Three\0"
@[c:'ImGui_ComboCallback']
fn combo_callback(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int) bool

// Implied popup_max_height_in_items = -1
@[c:'ImGui_ComboCallbackEx']
fn combo_callback_ex(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int, popup_max_height_in_items int) bool

// Widgets: Drag Sliders
// - CTRL+Click on any drag box to turn them into an input box. Manually input values aren't clamped by default and can go off-bounds. Use SliderFlags_AlwaysClamp to always clamp.
// - For all the Float2/Float3/Float4/Int2/Int3/Int4 versions of every function, note that a 'float v[X]' function argument is the same as 'float* v',
//   the array syntax is just a way to document the number of elements that are expected to be accessible. You can pass address of your first element out of a contiguous set, e.g. &myvector.x
// - Adjust format string to decorate the value with a prefix, a suffix, or adapt the editing and display precision e.g. "%.3f" -> 1.234; "%5.2f secs" -> 01.23 secs; "Biscuit: %.0f" -> Biscuit: 1; etc.
// - Format string may also be set to NULL or use the default format ("%f" or "%d").
// - Speed are per-pixel of mouse movement (v_speed=0.2f: mouse needs to move by 5 pixels to increase value by 1). For keyboard/gamepad navigation, minimum speed is Max(v_speed, minimum_step_at_given_precision).
// - Use v_min < v_max to clamp edits to given limits. Note that CTRL+Click manual input can override those limits if SliderFlags_AlwaysClamp is not used.
// - Use v_max = FLT_MAX / INT_MAX etc to avoid clamping to a maximum, same with v_min = -FLT_MAX / INT_MIN to avoid clamping to a minimum.
// - We use the same sets of flags for DragXXX() and SliderXXX() functions as the features are the same and it makes it easier to swap them.
// - Legacy: Pre-1.78 there are DragXXX() function signatures that take a final `float power=1.0f' argument instead of the  SliderFlags flags=0' argument.
//   If you get a warning converting a float to SliderFlags, read https://github.com/ocornut/imgui/issues/3361
@[c:'ImGui_DragFloat']
fn drag_float(label &i8, v &f32) bool

// Implied v_speed = 1.0f, v_min = 0.0f, v_max = 0.0f, format = "%.3f", flags = 0
@[c:'ImGui_DragFloatEx']
fn drag_float_ex(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

// If v_min >= v_max we have no bound
@[c:'ImGui_DragFloat2']
fn drag_float2(label &i8, v &f32) bool

// Implied v_speed = 1.0f, v_min = 0.0f, v_max = 0.0f, format = "%.3f", flags = 0
@[c:'ImGui_DragFloat2Ex']
fn drag_float2_ex(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragFloat3']
fn drag_float3(label &i8, v &f32) bool

// Implied v_speed = 1.0f, v_min = 0.0f, v_max = 0.0f, format = "%.3f", flags = 0
@[c:'ImGui_DragFloat3Ex']
fn drag_float3_ex(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragFloat4']
fn drag_float4(label &i8, v &f32) bool

// Implied v_speed = 1.0f, v_min = 0.0f, v_max = 0.0f, format = "%.3f", flags = 0
@[c:'ImGui_DragFloat4Ex']
fn drag_float4_ex(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragFloatRange2']
fn drag_float_range2(label &i8, v_current_min &f32, v_current_max &f32) bool

// Implied v_speed = 1.0f, v_min = 0.0f, v_max = 0.0f, format = "%.3f", format_max = NULL, flags = 0
@[c:'ImGui_DragFloatRange2Ex']
fn drag_float_range2_ex(label &i8, v_current_min &f32, v_current_max &f32, v_speed f32, v_min f32, v_max f32, format &i8, format_max &i8, flags SliderFlags) bool

@[c:'ImGui_DragInt']
fn drag_int(label &i8, v &int) bool

// Implied v_speed = 1.0f, v_min = 0, v_max = 0, format = "%d", flags = 0
@[c:'ImGui_DragIntEx']
fn drag_int_ex(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

// If v_min >= v_max we have no bound
@[c:'ImGui_DragInt2']
fn drag_int2(label &i8, v &int) bool

// Implied v_speed = 1.0f, v_min = 0, v_max = 0, format = "%d", flags = 0
@[c:'ImGui_DragInt2Ex']
fn drag_int2_ex(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragInt3']
fn drag_int3(label &i8, v &int) bool

// Implied v_speed = 1.0f, v_min = 0, v_max = 0, format = "%d", flags = 0
@[c:'ImGui_DragInt3Ex']
fn drag_int3_ex(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragInt4']
fn drag_int4(label &i8, v &int) bool

// Implied v_speed = 1.0f, v_min = 0, v_max = 0, format = "%d", flags = 0
@[c:'ImGui_DragInt4Ex']
fn drag_int4_ex(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragIntRange2']
fn drag_int_range2(label &i8, v_current_min &int, v_current_max &int) bool

// Implied v_speed = 1.0f, v_min = 0, v_max = 0, format = "%d", format_max = NULL, flags = 0
@[c:'ImGui_DragIntRange2Ex']
fn drag_int_range2_ex(label &i8, v_current_min &int, v_current_max &int, v_speed f32, v_min int, v_max int, format &i8, format_max &i8, flags SliderFlags) bool

@[c:'ImGui_DragScalar']
fn drag_scalar(label &i8, data_type DataType, p_data voidptr) bool

// Implied v_speed = 1.0f, p_min = NULL, p_max = NULL, format = NULL, flags = 0
@[c:'ImGui_DragScalarEx']
fn drag_scalar_ex(label &i8, data_type DataType, p_data voidptr, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c:'ImGui_DragScalarN']
fn drag_scalar_n(label &i8, data_type DataType, p_data voidptr, components int) bool

// Implied v_speed = 1.0f, p_min = NULL, p_max = NULL, format = NULL, flags = 0
@[c:'ImGui_DragScalarNEx']
fn drag_scalar_ne_x(label &i8, data_type DataType, p_data voidptr, components int, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

// Widgets: Regular Sliders
// - CTRL+Click on any slider to turn them into an input box. Manually input values aren't clamped by default and can go off-bounds. Use SliderFlags_AlwaysClamp to always clamp.
// - Adjust format string to decorate the value with a prefix, a suffix, or adapt the editing and display precision e.g. "%.3f" -> 1.234; "%5.2f secs" -> 01.23 secs; "Biscuit: %.0f" -> Biscuit: 1; etc.
// - Format string may also be set to NULL or use the default format ("%f" or "%d").
// - Legacy: Pre-1.78 there are SliderXXX() function signatures that take a final `float power=1.0f' argument instead of the  SliderFlags flags=0' argument.
//   If you get a warning converting a float to SliderFlags, read https://github.com/ocornut/imgui/issues/3361
@[c:'ImGui_SliderFloat']
fn slider_float(label &i8, v &f32, v_min f32, v_max f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_SliderFloatEx']
fn slider_float_ex(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

// adjust format to decorate the value with a prefix or a suffix for in-slider labels or unit display.
@[c:'ImGui_SliderFloat2']
fn slider_float2(label &i8, v &f32, v_min f32, v_max f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_SliderFloat2Ex']
fn slider_float2_ex(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderFloat3']
fn slider_float3(label &i8, v &f32, v_min f32, v_max f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_SliderFloat3Ex']
fn slider_float3_ex(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderFloat4']
fn slider_float4(label &i8, v &f32, v_min f32, v_max f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_SliderFloat4Ex']
fn slider_float4_ex(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderAngle']
fn slider_angle(label &i8, v_rad &f32) bool

// Implied v_degrees_min = -360.0f, v_degrees_max = +360.0f, format = "%.0f deg", flags = 0
@[c:'ImGui_SliderAngleEx']
fn slider_angle_ex(label &i8, v_rad &f32, v_degrees_min f32, v_degrees_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderInt']
fn slider_int(label &i8, v &int, v_min int, v_max int) bool

// Implied format = "%d", flags = 0
@[c:'ImGui_SliderIntEx']
fn slider_int_ex(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderInt2']
fn slider_int2(label &i8, v &int, v_min int, v_max int) bool

// Implied format = "%d", flags = 0
@[c:'ImGui_SliderInt2Ex']
fn slider_int2_ex(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderInt3']
fn slider_int3(label &i8, v &int, v_min int, v_max int) bool

// Implied format = "%d", flags = 0
@[c:'ImGui_SliderInt3Ex']
fn slider_int3_ex(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderInt4']
fn slider_int4(label &i8, v &int, v_min int, v_max int) bool

// Implied format = "%d", flags = 0
@[c:'ImGui_SliderInt4Ex']
fn slider_int4_ex(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderScalar']
fn slider_scalar(label &i8, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr) bool

// Implied format = NULL, flags = 0
@[c:'ImGui_SliderScalarEx']
fn slider_scalar_ex(label &i8, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c:'ImGui_SliderScalarN']
fn slider_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, p_min voidptr, p_max voidptr) bool

// Implied format = NULL, flags = 0
@[c:'ImGui_SliderScalarNEx']
fn slider_scalar_ne_x(label &i8, data_type DataType, p_data voidptr, components int, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c:'ImGui_VSliderFloat']
fn vs_lider_float(label &i8, size ImVec2, v &f32, v_min f32, v_max f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_VSliderFloatEx']
fn vs_lider_float_ex(label &i8, size ImVec2, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c:'ImGui_VSliderInt']
fn vs_lider_int(label &i8, size ImVec2, v &int, v_min int, v_max int) bool

// Implied format = "%d", flags = 0
@[c:'ImGui_VSliderIntEx']
fn vs_lider_int_ex(label &i8, size ImVec2, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c:'ImGui_VSliderScalar']
fn vs_lider_scalar(label &i8, size ImVec2, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr) bool

// Implied format = NULL, flags = 0
@[c:'ImGui_VSliderScalarEx']
fn vs_lider_scalar_ex(label &i8, size ImVec2, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

// Widgets: Input with Keyboard
// - If you want to use InputText() with std::string or any custom dynamic string type, see misc/cpp/imgui_stdlib.h and comments in imgui_demo.cpp.
// - Most of the InputTextFlags flags are only useful for InputText() and not for InputFloatX, InputIntX, InputDouble etc.
@[c:'ImGui_InputText']
fn input_text(label &i8, buf &i8, buf_size usize, flags InputTextFlags) bool

// Implied callback = NULL, user_data = NULL
@[c:'ImGui_InputTextEx']
fn input_text_ex(label &i8, buf &i8, buf_size usize, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c:'ImGui_InputTextMultiline']
fn input_text_multiline(label &i8, buf &i8, buf_size usize) bool

// Implied size = ImVec2(0, 0), flags = 0, callback = NULL, user_data = NULL
@[c:'ImGui_InputTextMultilineEx']
fn input_text_multiline_ex(label &i8, buf &i8, buf_size usize, size ImVec2, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c:'ImGui_InputTextWithHint']
fn input_text_with_hint(label &i8, hint &i8, buf &i8, buf_size usize, flags InputTextFlags) bool

// Implied callback = NULL, user_data = NULL
@[c:'ImGui_InputTextWithHintEx']
fn input_text_with_hint_ex(label &i8, hint &i8, buf &i8, buf_size usize, flags InputTextFlags, callback C.ImGuiInputTextCallback, user_data voidptr) bool

@[c:'ImGui_InputFloat']
fn input_float(label &i8, v &f32) bool

// Implied step = 0.0f, step_fast = 0.0f, format = "%.3f", flags = 0
@[c:'ImGui_InputFloatEx']
fn input_float_ex(label &i8, v &f32, step f32, step_fast f32, format &i8, flags InputTextFlags) bool

@[c:'ImGui_InputFloat2']
fn input_float2(label &i8, v &f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_InputFloat2Ex']
fn input_float2_ex(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c:'ImGui_InputFloat3']
fn input_float3(label &i8, v &f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_InputFloat3Ex']
fn input_float3_ex(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c:'ImGui_InputFloat4']
fn input_float4(label &i8, v &f32) bool

// Implied format = "%.3f", flags = 0
@[c:'ImGui_InputFloat4Ex']
fn input_float4_ex(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c:'ImGui_InputInt']
fn input_int(label &i8, v &int) bool

// Implied step = 1, step_fast = 100, flags = 0
@[c:'ImGui_InputIntEx']
fn input_int_ex(label &i8, v &int, step int, step_fast int, flags InputTextFlags) bool

@[c:'ImGui_InputInt2']
fn input_int2(label &i8, v &int, flags InputTextFlags) bool

@[c:'ImGui_InputInt3']
fn input_int3(label &i8, v &int, flags InputTextFlags) bool

@[c:'ImGui_InputInt4']
fn input_int4(label &i8, v &int, flags InputTextFlags) bool

@[c:'ImGui_InputDouble']
fn input_double(label &i8, v &f64) bool

// Implied step = 0.0, step_fast = 0.0, format = "%.6f", flags = 0
@[c:'ImGui_InputDoubleEx']
fn input_double_ex(label &i8, v &f64, step f64, step_fast f64, format &i8, flags InputTextFlags) bool

@[c:'ImGui_InputScalar']
fn input_scalar(label &i8, data_type DataType, p_data voidptr) bool

// Implied p_step = NULL, p_step_fast = NULL, format = NULL, flags = 0
@[c:'ImGui_InputScalarEx']
fn input_scalar_ex(label &i8, data_type DataType, p_data voidptr, p_step voidptr, p_step_fast voidptr, format &i8, flags InputTextFlags) bool

@[c:'ImGui_InputScalarN']
fn input_scalar_n(label &i8, data_type DataType, p_data voidptr, components int) bool

// Implied p_step = NULL, p_step_fast = NULL, format = NULL, flags = 0
@[c:'ImGui_InputScalarNEx']
fn input_scalar_ne_x(label &i8, data_type DataType, p_data voidptr, components int, p_step voidptr, p_step_fast voidptr, format &i8, flags InputTextFlags) bool

// Widgets: Color Editor/Picker (tip: the ColorEdit* functions have a little color square that can be left-clicked to open a picker, and right-clicked to open an option menu.)
// - Note that in C++ a 'float v[X]' function argument is the _same_ as 'float* v', the array syntax is just a way to document the number of elements that are expected to be accessible.
// - You can pass the address of a first float element out of a contiguous structure, e.g. &myvector.x
@[c:'ImGui_ColorEdit3']
fn color_edit3(label &i8, col &f32, flags ColorEditFlags) bool

@[c:'ImGui_ColorEdit4']
fn color_edit4(label &i8, col &f32, flags ColorEditFlags) bool

@[c:'ImGui_ColorPicker3']
fn color_picker3(label &i8, col &f32, flags ColorEditFlags) bool

@[c:'ImGui_ColorPicker4']
fn color_picker4(label &i8, col &f32, flags ColorEditFlags, ref_col &f32) bool

@[c:'ImGui_ColorButton']
fn color_button(desc_id &i8, col C.ImVec4, flags ColorEditFlags) bool

// Implied size = ImVec2(0, 0)
@[c:'ImGui_ColorButtonEx']
fn color_button_ex(desc_id &i8, col C.ImVec4, flags ColorEditFlags, size ImVec2) bool

// display a color square/button, hover for details, return true when pressed.
@[c:'ImGui_SetColorEditOptions']
fn set_color_edit_options(flags ColorEditFlags)

// initialize current options (generally on application startup) if you want to select a default format, picker type, etc. User will be able to change many settings, unless you pass the _NoOptions flag to your calls.
// Widgets: Trees
// - TreeNode functions return true when the node is open, in which case you need to also call TreePop() when you are finished displaying the tree node contents.
@[c:'ImGui_TreeNode']
fn tree_node(label &i8) bool

@[c2v_variadic]
@[c:'ImGui_TreeNodeStr']
fn tree_node_str(str_id &i8, fmt &i8) bool

// helper variation to easily decorelate the id from the displayed string. Read the FAQ about why and how to use ID. to align arbitrary text at the same level as a TreeNode() you can use Bullet().
@[c2v_variadic]
@[c:'ImGui_TreeNodePtr']
fn tree_node_ptr(ptr_id voidptr, fmt &i8) bool

// "
@[c:'ImGui_TreeNodeV']
fn tree_node_v(str_id &i8, fmt &i8, args C.va_list) bool

@[c:'ImGui_TreeNodeVPtr']
fn tree_node_vp_tr(ptr_id voidptr, fmt &i8, args C.va_list) bool

@[c:'ImGui_TreeNodeEx']
fn tree_node_ex(label &i8, flags TreeNodeFlags) bool

@[c2v_variadic]
@[c:'ImGui_TreeNodeExStr']
fn tree_node_ex_str(str_id &i8, flags TreeNodeFlags, fmt &i8) bool

@[c2v_variadic]
@[c:'ImGui_TreeNodeExPtr']
fn tree_node_ex_ptr(ptr_id voidptr, flags TreeNodeFlags, fmt &i8) bool

@[c:'ImGui_TreeNodeExV']
fn tree_node_ex_v(str_id &i8, flags TreeNodeFlags, fmt &i8, args C.va_list) bool

@[c:'ImGui_TreeNodeExVPtr']
fn tree_node_ex_vp_tr(ptr_id voidptr, flags TreeNodeFlags, fmt &i8, args C.va_list) bool

@[c:'ImGui_TreePush']
fn tree_push(str_id &i8)

// ~ Indent()+PushID(). Already called by TreeNode() when returning true, but you can call TreePush/TreePop yourself if desired.
@[c:'ImGui_TreePushPtr']
fn tree_push_ptr(ptr_id voidptr)

// "
@[c:'ImGui_TreePop']
fn tree_pop()

// ~ Unindent()+PopID()
@[c:'ImGui_GetTreeNodeToLabelSpacing']
fn get_tree_node_to_label_spacing() f32

// horizontal distance preceding label when using TreeNode*() or Bullet() == (g.FontSize + style.FramePadding.x*2) for a regular unframed TreeNode
@[c:'ImGui_CollapsingHeader']
fn collapsing_header(label &i8, flags TreeNodeFlags) bool

// if returning 'true' the header is open. doesn't indent nor push on ID stack. user doesn't have to call TreePop().
@[c:'ImGui_CollapsingHeaderBoolPtr']
fn collapsing_header_bool_ptr(label &i8, p_visible &bool, flags TreeNodeFlags) bool

// when 'p_visible != NULL': if '*p_visible==true' display an additional small close button on upper right of the header which will set the bool to false when clicked, if '*p_visible==false' don't display the header.
@[c:'ImGui_SetNextItemOpen']
fn set_next_item_open(is_open bool, cond Cond)

// set next TreeNode/CollapsingHeader open state.
@[c:'ImGui_SetNextItemStorageID']
fn set_next_item_storage_id(storage_id ID)

// set id to use for open/close storage (default to same as item id).
// Widgets: Selectables
// - A selectable highlights when hovered, and can display another color when selected.
// - Neighbors selectable extend their highlight bounds in order to leave no gap between them. This is so a series of selected Selectable appear contiguous.
@[c:'ImGui_Selectable']
fn selectable(label &i8) bool

// Implied selected = false, flags = 0, size = ImVec2(0, 0)
@[c:'ImGui_SelectableEx']
fn selectable_ex(label &i8, selected bool, flags SelectableFlags, size ImVec2) bool

// "bool selected" carry the selection state (read-only). Selectable() is clicked is returns true so you can modify your selection state. size.x==0.0: use remaining width, size.x>0.0: specify width. size.y==0.0: use label height, size.y>0.0: specify height
@[c:'ImGui_SelectableBoolPtr']
fn selectable_bool_ptr(label &i8, p_selected &bool, flags SelectableFlags) bool

// Implied size = ImVec2(0, 0)
@[c:'ImGui_SelectableBoolPtrEx']
fn selectable_bool_ptr_ex(label &i8, p_selected &bool, flags SelectableFlags, size ImVec2) bool

// "bool* p_selected" point to the selection state (read-write), as a convenient helper.
// Multi-selection system for Selectable(), Checkbox(), TreeNode() functions [BETA]
// - This enables standard multi-selection/range-selection idioms (CTRL+Mouse/Keyboard, SHIFT+Mouse/Keyboard, etc.) in a way that also allow a clipper to be used.
// - SelectionUserData is often used to store your item index within the current view (but may store something else).
// - Read comments near ImGuiMultiSelectIO for instructions/details and see 'Demo->Widgets->Selection State & Multi-Select' for demo.
// - TreeNode() is technically supported but... using this correctly is more complicated. You need some sort of linear/random access to your tree,
//   which is suited to advanced trees setups already implementing filters and clipper. We will work simplifying the current demo.
// - 'selection_size' and 'items_count' parameters are optional and used by a few features. If they are costly for you to compute, you may avoid them.
@[c:'ImGui_BeginMultiSelect']
fn begin_multi_select(flags MultiSelectFlags) &ImGuiMultiSelectIO

// Implied selection_size = -1, items_count = -1
@[c:'ImGui_BeginMultiSelectEx']
fn begin_multi_select_ex(flags MultiSelectFlags, selection_size int, items_count int) &ImGuiMultiSelectIO

@[c:'ImGui_EndMultiSelect']
fn end_multi_select() &ImGuiMultiSelectIO

@[c:'ImGui_SetNextItemSelectionUserData']
fn set_next_item_selection_user_data(selection_user_data SelectionUserData)

@[c:'ImGui_IsItemToggledSelection']
fn is_item_toggled_selection() bool

// Was the last item selection state toggled? Useful if you need the per-item information _before_ reaching EndMultiSelect(). We only returns toggle _event_ in order to handle clipping correctly.
// Widgets: List Boxes
// - This is essentially a thin wrapper to using BeginChild/EndChild with the ChildFlags_FrameStyle flag for stylistic changes + displaying a label.
// - If you don't need a label you can probably simply use BeginChild() with the ChildFlags_FrameStyle flag for the same result.
// - You can submit contents and manage your selection state however you want it, by creating e.g. Selectable() or any other items.
// - The simplified/old ListBox() api are helpers over BeginListBox()/EndListBox() which are kept available for convenience purpose. This is analoguous to how Combos are created.
// - Choose frame width:   size.x > 0.0f: custom  /  size.x < 0.0f or -FLT_MIN: right-align   /  size.x = 0.0f (default): use current ItemWidth
// - Choose frame height:  size.y > 0.0f: custom  /  size.y < 0.0f or -FLT_MIN: bottom-align  /  size.y = 0.0f (default): arbitrary default height which can fit ~7 items
@[c:'ImGui_BeginListBox']
fn begin_list_box(label &i8, size ImVec2) bool

// open a framed scrolling region
@[c:'ImGui_EndListBox']
fn end_list_box()

// only call EndListBox() if BeginListBox() returned true!
@[c:'ImGui_ListBox']
fn list_box(label &i8, current_item &int, items &&u8, items_count int, height_in_items int) bool

@[c:'ImGui_ListBoxCallback']
fn list_box_callback(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int) bool

// Implied height_in_items = -1
@[c:'ImGui_ListBoxCallbackEx']
fn list_box_callback_ex(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int, height_in_items int) bool

// Widgets: Data Plotting
// - Consider using ImPlot (https://github.com/epezent/implot) which is much better!
@[c:'ImGui_PlotLines']
fn plot_lines(label &i8, values &f32, values_count int)

// Implied values_offset = 0, overlay_text = NULL, scale_min = FLT_MAX, scale_max = FLT_MAX, graph_size = ImVec2(0, 0), stride = sizeof(float)
@[c:'ImGui_PlotLinesEx']
fn plot_lines_ex(label &i8, values &f32, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2, stride int)

@[c:'ImGui_PlotLinesCallback']
fn plot_lines_callback(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int)

// Implied values_offset = 0, overlay_text = NULL, scale_min = FLT_MAX, scale_max = FLT_MAX, graph_size = ImVec2(0, 0)
@[c:'ImGui_PlotLinesCallbackEx']
fn plot_lines_callback_ex(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2)

@[c:'ImGui_PlotHistogram']
fn plot_histogram(label &i8, values &f32, values_count int)

// Implied values_offset = 0, overlay_text = NULL, scale_min = FLT_MAX, scale_max = FLT_MAX, graph_size = ImVec2(0, 0), stride = sizeof(float)
@[c:'ImGui_PlotHistogramEx']
fn plot_histogram_ex(label &i8, values &f32, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2, stride int)

@[c:'ImGui_PlotHistogramCallback']
fn plot_histogram_callback(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int)

// Implied values_offset = 0, overlay_text = NULL, scale_min = FLT_MAX, scale_max = FLT_MAX, graph_size = ImVec2(0, 0)
@[c:'ImGui_PlotHistogramCallbackEx']
fn plot_histogram_callback_ex(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2)

// Widgets: Menus
// - Use BeginMenuBar() on a window WindowFlags_MenuBar to append to its menu bar.
// - Use BeginMainMenuBar() to create a menu bar at the top of the screen and append to it.
// - Use BeginMenu() to create a menu. You can call BeginMenu() multiple time with the same identifier to append more items to it.
// - Not that MenuItem() keyboardshortcuts are displayed as a convenience but _not processed_ by Dear ImGui at the moment.
@[c:'ImGui_BeginMenuBar']
fn begin_menu_bar() bool

// append to menu-bar of current window (requires WindowFlags_MenuBar flag set on parent window).
@[c:'ImGui_EndMenuBar']
fn end_menu_bar()

// only call EndMenuBar() if BeginMenuBar() returns true!
@[c:'ImGui_BeginMainMenuBar']
fn begin_main_menu_bar() bool

// create and append to a full screen menu-bar.
@[c:'ImGui_EndMainMenuBar']
fn end_main_menu_bar()

// only call EndMainMenuBar() if BeginMainMenuBar() returns true!
@[c:'ImGui_BeginMenu']
fn begin_menu(label &i8) bool

// Implied enabled = true
@[c:'ImGui_BeginMenuEx']
fn begin_menu_ex(label &i8, enabled bool) bool

// create a sub-menu entry. only call EndMenu() if this returns true!
@[c:'ImGui_EndMenu']
fn end_menu()

// only call EndMenu() if BeginMenu() returns true!
@[c:'ImGui_MenuItem']
fn menu_item(label &i8) bool

// Implied shortcut = NULL, selected = false, enabled = true
@[c:'ImGui_MenuItemEx']
fn menu_item_ex(label &i8, shortcut &i8, selected bool, enabled bool) bool

// return true when activated.
@[c:'ImGui_MenuItemBoolPtr']
fn menu_item_bool_ptr(label &i8, shortcut &i8, p_selected &bool, enabled bool) bool

// return true when activated + toggle (*p_selected) if p_selected != NULL
// Tooltips
// - Tooltips are windows following the mouse. They do not take focus away.
// - A tooltip window can contain items of any types.
// - SetTooltip() is more or less a shortcut for the 'if (BeginTooltip()) { Text(...); EndTooltip(); }' idiom (with a subtlety that it discard any previously submitted tooltip)
@[c:'ImGui_BeginTooltip']
fn begin_tooltip() bool

// begin/append a tooltip window.
@[c:'ImGui_EndTooltip']
fn end_tooltip()

// only call EndTooltip() if BeginTooltip()/BeginItemTooltip() returns true!
@[c2v_variadic]
@[c:'ImGui_SetTooltip']
fn set_tooltip(fmt &i8)

// set a text-only tooltip. Often used after a ImGui::IsItemHovered() check. Override any previous call to SetTooltip().
@[c:'ImGui_SetTooltipV']
fn set_tooltip_v(fmt &i8, args C.va_list)

// Tooltips: helpers for showing a tooltip when hovering an item
// - BeginItemTooltip() is a shortcut for the 'if (IsItemHovered HoveredFlags_ForTooltip) && BeginTooltip())' idiom.
// - SetItemTooltip() is a shortcut for the 'if (IsItemHovered HoveredFlags_ForTooltip)) { SetTooltip(...); }' idiom.
// - Where 'ImGuiHoveredFlags_ForTooltip' itself is a shortcut to use 'style.HoverFlagsForTooltipMouse' or 'style.HoverFlagsForTooltipNav' depending on active input type. For mouse it defaults to 'ImGuiHoveredFlags_Stationary | HoveredFlags_DelayShort'.
@[c:'ImGui_BeginItemTooltip']
fn begin_item_tooltip() bool

// begin/append a tooltip window if preceding item was hovered.
@[c2v_variadic]
@[c:'ImGui_SetItemTooltip']
fn set_item_tooltip(fmt &i8)

// set a text-only tooltip if preceding item was hovered. override any previous call to SetTooltip().
@[c:'ImGui_SetItemTooltipV']
fn set_item_tooltip_v(fmt &i8, args C.va_list)

// Popups, Modals
//  - They block normal mouse hovering detection (and therefore most mouse interactions) behind them.
//  - If not modal: they can be closed by clicking anywhere outside them, or by pressing ESCAPE.
//  - Their visibility state (~bool) is held internally instead of being held by the programmer as we are used to with regular Begin*() calls.
//  - The 3 properties above are related: we need to retain popup visibility state in the library because popups may be closed as any time.
//  - You can bypass the hovering restriction by using HoveredFlags_AllowWhenBlockedByPopup when calling IsItemHovered() or IsWindowHovered().
//  - IMPORTANT: Popup identifiers are relative to the current ID stack, so OpenPopup and BeginPopup generally needs to be at the same level of the stack.
//    This is sometimes leading to confusing mistakes. May rework this in the future.
//  - BeginPopup(): query popup state, if open start appending into the window. Call EndPopup() afterwards if returned true. WindowFlags are forwarded to the window.
//  - BeginPopupModal(): block every interaction behind the window, cannot be closed by user, add a dimming background, has a title bar.
@[c:'ImGui_BeginPopup']
fn begin_popup(str_id &i8, flags WindowFlags) bool

// return true if the popup is open, and you can start outputting to it.
@[c:'ImGui_BeginPopupModal']
fn begin_popup_modal(name &i8, p_open &bool, flags WindowFlags) bool

// return true if the modal is open, and you can start outputting to it.
@[c:'ImGui_EndPopup']
fn end_popup()

// only call EndPopup() if BeginPopupXXX() returns true!
// Popups: open/close functions
//  - OpenPopup(): set popup state to open. PopupFlags are available for opening options.
//  - If not modal: they can be closed by clicking anywhere outside them, or by pressing ESCAPE.
//  - CloseCurrentPopup(): use inside the BeginPopup()/EndPopup() scope to close manually.
//  - CloseCurrentPopup() is called by default by Selectable()/MenuItem() when activated (FIXME: need some options).
//  - Use PopupFlags_NoOpenOverExistingPopup to avoid opening a popup if there's already one at the same level. This is equivalent to e.g. testing for !IsAnyPopupOpen() prior to OpenPopup().
//  - Use IsWindowAppearing() after BeginPopup() to tell if a window just opened.
//  - IMPORTANT: Notice that for OpenPopupOnItemClick() we exceptionally default flags to 1 (== PopupFlags_MouseButtonRight) for backward compatibility with older API taking 'int mouse_button = 1' parameter
@[c:'ImGui_OpenPopup']
fn open_popup(str_id &i8, popup_flags PopupFlags)

// call to mark popup as open (don't call every frame!).
@[c:'ImGui_OpenPopupID']
fn open_popup_id(id ID, popup_flags PopupFlags)

// id overload to facilitate calling from nested stacks
@[c:'ImGui_OpenPopupOnItemClick']
fn open_popup_on_item_click(str_id &i8, popup_flags PopupFlags)

// helper to open popup when clicked on last item. Default to PopupFlags_MouseButtonRight == 1. (note: actually triggers on the mouse _released_ event to be consistent with popup behaviors)
@[c:'ImGui_CloseCurrentPopup']
fn close_current_popup()

// manually close the popup we have begin-ed into.
// Popups: open+begin combined functions helpers
//  - Helpers to do OpenPopup+BeginPopup where the Open action is triggered by e.g. hovering an item and right-clicking.
//  - They are convenient to easily create context menus, hence the name.
//  - IMPORTANT: Notice that BeginPopupContextXXX takes PopupFlags just like OpenPopup() and unlike BeginPopup(). For full consistency, we may add WindowFlags to the BeginPopupContextXXX functions in the future.
//  - IMPORTANT: Notice that we exceptionally default their flags to 1 (== PopupFlags_MouseButtonRight) for backward compatibility with older API taking 'int mouse_button = 1' parameter, so if you add other flags remember to re-add the PopupFlags_MouseButtonRight.
@[c:'ImGui_BeginPopupContextItem']
fn begin_popup_context_item() bool

// Implied str_id = NULL, popup_flags = 1
@[c:'ImGui_BeginPopupContextItemEx']
fn begin_popup_context_item_ex(str_id &i8, popup_flags PopupFlags) bool

// open+begin popup when clicked on last item. Use str_id==NULL to associate the popup to previous item. If you want to use that on a non-interactive item such as Text() you need to pass in an explicit ID here. read comments in .cpp!
@[c:'ImGui_BeginPopupContextWindow']
fn begin_popup_context_window() bool

// Implied str_id = NULL, popup_flags = 1
@[c:'ImGui_BeginPopupContextWindowEx']
fn begin_popup_context_window_ex(str_id &i8, popup_flags PopupFlags) bool

// open+begin popup when clicked on current window.
@[c:'ImGui_BeginPopupContextVoid']
fn begin_popup_context_void() bool

// Implied str_id = NULL, popup_flags = 1
@[c:'ImGui_BeginPopupContextVoidEx']
fn begin_popup_context_void_ex(str_id &i8, popup_flags PopupFlags) bool

// open+begin popup when clicked in void (where there are no windows).
// Popups: query functions
//  - IsPopupOpen(): return true if the popup is open at the current BeginPopup() level of the popup stack.
//  - IsPopupOpen() with PopupFlags_AnyPopupId: return true if any popup is open at the current BeginPopup() level of the popup stack.
//  - IsPopupOpen() with PopupFlags_AnyPopupId + PopupFlags_AnyPopupLevel: return true if any popup is open.
@[c:'ImGui_IsPopupOpen']
fn is_popup_open(str_id &i8, flags PopupFlags) bool

// return true if the popup is open.
// Tables
// - Full-featured replacement for old Columns API.
// - See Demo->Tables for demo code. See top of imgui_tables.cpp for general commentary.
// - See TableFlags_ and TableColumnFlags_ enums for a description of available flags.
// The typical call flow is:
// - 1. Call BeginTable(), early out if returning false.
// - 2. Optionally call TableSetupColumn() to submit column name/flags/defaults.
// - 3. Optionally call TableSetupScrollFreeze() to request scroll freezing of columns/rows.
// - 4. Optionally call TableHeadersRow() to submit a header row. Names are pulled from TableSetupColumn() data.
// - 5. Populate contents:
//    - In most situations you can use TableNextRow() + TableSetColumnIndex(N) to start appending into a column.
//    - If you are using tables as a sort of grid, where every column is holding the same type of contents,
//      you may prefer using TableNextColumn() instead of TableNextRow() + TableSetColumnIndex().
//      TableNextColumn() will automatically wrap-around into the next row if needed.
//    - IMPORTANT: Comparatively to the old Columns() API, we need to call TableNextColumn() for the first column!
//    - Summary of possible call flow:
//        - TableNextRow() -> TableSetColumnIndex(0) -> Text("Hello 0") -> TableSetColumnIndex(1) -> Text("Hello 1")  // OK
//        - TableNextRow() -> TableNextColumn()      -> Text("Hello 0") -> TableNextColumn()      -> Text("Hello 1")  // OK
//        -                   TableNextColumn()      -> Text("Hello 0") -> TableNextColumn()      -> Text("Hello 1")  // OK: TableNextColumn() automatically gets to next row!
//        - TableNextRow()                           -> Text("Hello 0")                                               // Not OK! Missing TableSetColumnIndex() or TableNextColumn()! Text will not appear!
// - 5. Call EndTable()
@[c:'ImGui_BeginTable']
fn begin_table(str_id &i8, columns int, flags TableFlags) bool

// Implied outer_size = ImVec2(0.0f, 0.0f), inner_width = 0.0f
@[c:'ImGui_BeginTableEx']
fn begin_table_ex(str_id &i8, columns int, flags TableFlags, outer_size ImVec2, inner_width f32) bool

@[c:'ImGui_EndTable']
fn end_table()

// only call EndTable() if BeginTable() returns true!
@[c:'ImGui_TableNextRow']
fn table_next_row()

// Implied row_flags = 0, min_row_height = 0.0f
@[c:'ImGui_TableNextRowEx']
fn table_next_row_ex(row_flags TableRowFlags, min_row_height f32)

// append into the first cell of a new row.
@[c:'ImGui_TableNextColumn']
fn table_next_column() bool

// append into the next column (or first column of next row if currently in last column). Return true when column is visible.
@[c:'ImGui_TableSetColumnIndex']
fn table_set_column_index(column_n int) bool

// append into the specified column. Return true when column is visible.
// Tables: Headers & Columns declaration
// - Use TableSetupColumn() to specify label, resizing policy, default width/weight, id, various other flags etc.
// - Use TableHeadersRow() to create a header row and automatically submit a TableHeader() for each column.
//   Headers are required to perform: reordering, sorting, and opening the context menu.
//   The context menu can also be made available in columns body using TableFlags_ContextMenuInBody.
// - You may manually submit headers using TableNextRow() + TableHeader() calls, but this is only useful in
//   some advanced use cases (e.g. adding custom widgets in header row).
// - Use TableSetupScrollFreeze() to lock columns/rows so they stay visible when scrolled.
@[c:'ImGui_TableSetupColumn']
fn table_setup_column(label &i8, flags TableColumnFlags)

// Implied init_width_or_weight = 0.0f, user_id = 0
@[c:'ImGui_TableSetupColumnEx']
fn table_setup_column_ex(label &i8, flags TableColumnFlags, init_width_or_weight f32, user_id ID)

@[c:'ImGui_TableSetupScrollFreeze']
fn table_setup_scroll_freeze(cols int, rows int)

// lock columns/rows so they stay visible when scrolled.
@[c:'ImGui_TableHeader']
fn table_header(label &i8)

// submit one header cell manually (rarely used)
@[c:'ImGui_TableHeadersRow']
fn table_headers_row()

// submit a row with headers cells based on data provided to TableSetupColumn() + submit context menu
@[c:'ImGui_TableAngledHeadersRow']
fn table_angled_headers_row()

// submit a row with angled headers for every column with the TableColumnFlags_AngledHeader flag. MUST BE FIRST ROW.
// Tables: Sorting & Miscellaneous functions
// - Sorting: call TableGetSortSpecs() to retrieve latest sort specs for the table. NULL when not sorting.
//   When 'sort_specs->SpecsDirty == true' you should sort your data. It will be true when sorting specs have
//   changed since last call, or the first time. Make sure to set 'SpecsDirty = false' after sorting,
//   else you may wastefully sort your data every frame!
// - Functions args 'int column_n' treat the default value of -1 as the same as passing the current column index.
@[c:'ImGui_TableGetSortSpecs']
fn table_get_sort_specs() &ImGuiTableSortSpecs

// get latest sort specs for the table (NULL if not sorting).  Lifetime: don't hold on this pointer over multiple frames or past any subsequent call to BeginTable().
@[c:'ImGui_TableGetColumnCount']
fn table_get_column_count() int

// return number of columns (value passed to BeginTable)
@[c:'ImGui_TableGetColumnIndex']
fn table_get_column_index() int

// return current column index.
@[c:'ImGui_TableGetRowIndex']
fn table_get_row_index() int

// return current row index.
@[c:'ImGui_TableGetColumnName']
fn table_get_column_name(column_n int) &i8

// return "" if column didn't have a name declared by TableSetupColumn(). Pass -1 to use current column.
@[c:'ImGui_TableGetColumnFlags']
fn table_get_column_flags(column_n int) TableColumnFlags

// return column flags so you can query their Enabled/Visible/Sorted/Hovered status flags. Pass -1 to use current column.
@[c:'ImGui_TableSetColumnEnabled']
fn table_set_column_enabled(column_n int, v bool)

// change user accessible enabled/disabled state of a column. Set to false to hide the column. User can use the context menu to change this themselves (right-click in headers, or right-click in columns body with TableFlags_ContextMenuInBody)
@[c:'ImGui_TableGetHoveredColumn']
fn table_get_hovered_column() int

// return hovered column. return -1 when table is not hovered. return columns_count if the unused space at the right of visible columns is hovered. Can also use (TableGetColumnFlags() & TableColumnFlags_IsHovered) instead.
@[c:'ImGui_TableSetBgColor']
fn table_set_bg_color(target TableBgTarget, color ImU32, column_n int)

// change the color of a cell, row, or column. See TableBgTarget_ flags for details.
// Legacy Columns API (prefer using Tables!)
// - You can also use SameLine(pos_x) to mimic simplified columns.
@[c:'ImGui_Columns']
fn columns()

// Implied count = 1, id = NULL, borders = true
@[c:'ImGui_ColumnsEx']
fn columns_ex(count int, id &i8, borders bool)

@[c:'ImGui_NextColumn']
fn next_column()

// next column, defaults to current row or next row if the current row is finished
@[c:'ImGui_GetColumnIndex']
fn get_column_index() int

// get current column index
@[c:'ImGui_GetColumnWidth']
fn get_column_width(column_index int) f32

// get column width (in pixels). pass -1 to use current column
@[c:'ImGui_SetColumnWidth']
fn set_column_width(column_index int, width f32)

// set column width (in pixels). pass -1 to use current column
@[c:'ImGui_GetColumnOffset']
fn get_column_offset(column_index int) f32

// get position of column line (in pixels, from the left side of the contents region). pass -1 to use current column, otherwise 0..GetColumnsCount() inclusive. column 0 is typically 0.0f
@[c:'ImGui_SetColumnOffset']
fn set_column_offset(column_index int, offset_x f32)

// set position of column line (in pixels, from the left side of the contents region). pass -1 to use current column
@[c:'ImGui_GetColumnsCount']
fn get_columns_count() int

// Tab Bars, Tabs
// - Note: Tabs are automatically created by the docking system (when in 'docking' branch). Use this to create tab bars/tabs yourself.
@[c:'ImGui_BeginTabBar']
fn begin_tab_bar(str_id &i8, flags TabBarFlags) bool

// create and append into a TabBar
@[c:'ImGui_EndTabBar']
fn end_tab_bar()

// only call EndTabBar() if BeginTabBar() returns true!
@[c:'ImGui_BeginTabItem']
fn begin_tab_item(label &i8, p_open &bool, flags TabItemFlags) bool

// create a Tab. Returns true if the Tab is selected.
@[c:'ImGui_EndTabItem']
fn end_tab_item()

// only call EndTabItem() if BeginTabItem() returns true!
@[c:'ImGui_TabItemButton']
fn tab_item_button(label &i8, flags TabItemFlags) bool

// create a Tab behaving like a button. return true when clicked. cannot be selected in the tab bar.
@[c:'ImGui_SetTabItemClosed']
fn set_tab_item_closed(tab_or_docked_window_label &i8)

// notify TabBar or Docking system of a closed tab/window ahead (useful to reduce visual flicker on reorderable tab bars). For tab-bar: call after BeginTabBar() and before Tab submissions. Otherwise call with a window name.
// Logging/Capture
// - All text output from the interface can be captured into tty/file/clipboard. By default, tree nodes are automatically opened during logging.
@[c:'ImGui_LogToTTY']
fn log_to_tty(auto_open_depth int)

// start logging to tty (stdout)
@[c:'ImGui_LogToFile']
fn log_to_file(auto_open_depth int, filename &i8)

// start logging to file
@[c:'ImGui_LogToClipboard']
fn log_to_clipboard(auto_open_depth int)

// start logging to OS clipboard
@[c:'ImGui_LogFinish']
fn log_finish()

// stop logging (close file, etc.)
@[c:'ImGui_LogButtons']
fn log_buttons()

// helper to display buttons for logging to tty/file/clipboard
@[c2v_variadic]
@[c:'ImGui_LogText']
fn log_text(fmt &i8)

// pass text data straight to log (without being displayed)
@[c:'ImGui_LogTextV']
fn log_text_v(fmt &i8, args C.va_list)

// Drag and Drop
// - On source items, call BeginDragDropSource(), if it returns true also call SetDragDropPayload() + EndDragDropSource().
// - On target candidates, call BeginDragDropTarget(), if it returns true also call AcceptDragDropPayload() + EndDragDropTarget().
// - If you stop calling BeginDragDropSource() the payload is preserved however it won't have a preview tooltip (we currently display a fallback "..." tooltip, see #1725)
// - An item can be both drag source and drop target.
@[c:'ImGui_BeginDragDropSource']
fn begin_drag_drop_source(flags DragDropFlags) bool

// call after submitting an item which may be dragged. when this return true, you can call SetDragDropPayload() + EndDragDropSource()
@[c:'ImGui_SetDragDropPayload']
fn set_drag_drop_payload(type_ &i8, data voidptr, sz usize, cond Cond) bool

// type is a user defined string of maximum 32 characters. Strings starting with '_' are reserved for dear imgui internal types. Data is copied and held by imgui. Return true when payload has been accepted.
@[c:'ImGui_EndDragDropSource']
fn end_drag_drop_source()

// only call EndDragDropSource() if BeginDragDropSource() returns true!
@[c:'ImGui_BeginDragDropTarget']
fn begin_drag_drop_target() bool

// call after submitting an item that may receive a payload. If this returns true, you can call AcceptDragDropPayload() + EndDragDropTarget()
@[c:'ImGui_AcceptDragDropPayload']
fn accept_drag_drop_payload(type_ &i8, flags DragDropFlags) &ImGuiPayload

// accept contents of a given type. If DragDropFlags_AcceptBeforeDelivery is set you can peek into the payload before the mouse button is released.
@[c:'ImGui_EndDragDropTarget']
fn end_drag_drop_target()

// only call EndDragDropTarget() if BeginDragDropTarget() returns true!
@[c:'ImGui_GetDragDropPayload']
fn get_drag_drop_payload() &ImGuiPayload

// peek directly into the current payload from anywhere. returns NULL when drag and drop is finished or inactive. use ImGuiPayload::IsDataType() to test for the payload type.
// Disabling [BETA API]
// - Disable all user interactions and dim items visuals (applying style.DisabledAlpha over current colors)
// - Those can be nested but it cannot be used to enable an already disabled section (a single BeginDisabled(true) in the stack is enough to keep everything disabled)
// - Tooltips windows by exception are opted out of disabling.
// - BeginDisabled(false)/EndDisabled() essentially does nothing but is provided to facilitate use of boolean expressions (as a micro-optimization: if you have tens of thousands of BeginDisabled(false)/EndDisabled() pairs, you might want to reformulate your code to avoid making those calls)
@[c:'ImGui_BeginDisabled']
fn begin_disabled(disabled bool)

@[c:'ImGui_EndDisabled']
fn end_disabled()

// Clipping
// - Mouse hovering is affected by ImGui::PushClipRect() calls, unlike direct calls to ImDrawList::PushClipRect() which are render only.
@[c:'ImGui_PushClipRect']
fn push_clip_rect(clip_rect_min ImVec2, clip_rect_max ImVec2, intersect_with_current_clip_rect bool)

@[c:'ImGui_PopClipRect']
fn pop_clip_rect()

// Focus, Activation
@[c:'ImGui_SetItemDefaultFocus']
fn set_item_default_focus()

// make last item the default focused item of a newly appearing window.
@[c:'ImGui_SetKeyboardFocusHere']
fn set_keyboard_focus_here()

// Implied offset = 0
@[c:'ImGui_SetKeyboardFocusHereEx']
fn set_keyboard_focus_here_ex(offset int)

// focus keyboard on the next widget. Use positive 'offset' to access sub components of a multiple component widget. Use -1 to access previous widget.
// Keyboard/Gamepad Navigation
@[c:'ImGui_SetNavCursorVisible']
fn set_nav_cursor_visible(visible bool)

// alter visibility of keyboard/gamepad cursor. by default: show when using an arrow key, hide when clicking with mouse.
// Overlapping mode
@[c:'ImGui_SetNextItemAllowOverlap']
fn set_next_item_allow_overlap()

// allow next item to be overlapped by a subsequent item. Useful with invisible buttons, selectable, treenode covering an area where subsequent items may need to be added. Note that both Selectable() and TreeNode() have dedicated flags doing this.
// Item/Widgets Utilities and Query Functions
// - Most of the functions are referring to the previous Item that has been submitted.
// - See Demo Window under "Widgets->Querying Status" for an interactive visualization of most of those functions.
@[c:'ImGui_IsItemHovered']
fn is_item_hovered(flags HoveredFlags) bool

// is the last item hovered? (and usable, aka not blocked by a popup, etc.). See HoveredFlags for more options.
@[c:'ImGui_IsItemActive']
fn is_item_active() bool

// is the last item active? (e.g. button being held, text field being edited. This will continuously return true while holding mouse button on an item. Items that don't interact will always return false)
@[c:'ImGui_IsItemFocused']
fn is_item_focused() bool

// is the last item focused for keyboard/gamepad navigation?
@[c:'ImGui_IsItemClicked']
fn is_item_clicked() bool

// Implied mouse_button = 0
@[c:'ImGui_IsItemClickedEx']
fn is_item_clicked_ex(mouse_button MouseButton) bool

// is the last item hovered and mouse clicked on? (**)  == IsMouseClicked(mouse_button) && IsItemHovered()Important. (**) this is NOT equivalent to the behavior of e.g. Button(). Read comments in function definition.
@[c:'ImGui_IsItemVisible']
fn is_item_visible() bool

// is the last item visible? (items may be out of sight because of clipping/scrolling)
@[c:'ImGui_IsItemEdited']
fn is_item_edited() bool

// did the last item modify its underlying value this frame? or was pressed? This is generally the same as the "bool" return value of many widgets.
@[c:'ImGui_IsItemActivated']
fn is_item_activated() bool

// was the last item just made active (item was previously inactive).
@[c:'ImGui_IsItemDeactivated']
fn is_item_deactivated() bool

// was the last item just made inactive (item was previously active). Useful for Undo/Redo patterns with widgets that require continuous editing.
@[c:'ImGui_IsItemDeactivatedAfterEdit']
fn is_item_deactivated_after_edit() bool

// was the last item just made inactive and made a value change when it was active? (e.g. Slider/Drag moved). Useful for Undo/Redo patterns with widgets that require continuous editing. Note that you may get false positives (some widgets such as Combo()/ListBox()/Selectable() will return true even when clicking an already selected item).
@[c:'ImGui_IsItemToggledOpen']
fn is_item_toggled_open() bool

// was the last item open state toggled? set by TreeNode().
@[c:'ImGui_IsAnyItemHovered']
fn is_any_item_hovered() bool

// is any item hovered?
@[c:'ImGui_IsAnyItemActive']
fn is_any_item_active() bool

// is any item active?
@[c:'ImGui_IsAnyItemFocused']
fn is_any_item_focused() bool

// is any item focused?
@[c:'ImGui_GetItemID']
fn get_item_id() ID

// get ID of last item (~~ often same ImGui::GetID(label) beforehand)
@[c:'ImGui_GetItemRectMin']
fn get_item_rect_min() ImVec2

// get upper-left bounding rectangle of the last item (screen space)
@[c:'ImGui_GetItemRectMax']
fn get_item_rect_max() ImVec2

// get lower-right bounding rectangle of the last item (screen space)
@[c:'ImGui_GetItemRectSize']
fn get_item_rect_size() ImVec2

// get size of last item
// Viewports
// - Currently represents the Platform Window created by the application which is hosting our Dear ImGui windows.
// - In 'docking' branch with multi-viewport enabled, we extend this concept to have multiple active viewports.
// - In the future we will extend this concept further to also represent Platform Monitor and support a "no main platform window" operation mode.
@[c:'ImGui_GetMainViewport']
fn get_main_viewport() &ImGuiViewport

// return primary/default viewport. This can never be NULL.
// Background/Foreground Draw Lists
@[c:'ImGui_GetBackgroundDrawList']
fn get_background_draw_list() &ImDrawList

// this draw list will be the first rendered one. Useful to quickly draw shapes/text behind dear imgui contents.
@[c:'ImGui_GetForegroundDrawList']
fn get_foreground_draw_list() &ImDrawList

// this draw list will be the last rendered one. Useful to quickly draw shapes/text over dear imgui contents.
// Miscellaneous Utilities
@[c:'ImGui_IsRectVisibleBySize']
fn is_rect_visible_by_size(size ImVec2) bool

// test if rectangle (of given size, starting from cursor position) is visible / not clipped.
@[c:'ImGui_IsRectVisible']
fn is_rect_visible(rect_min ImVec2, rect_max ImVec2) bool

// test if rectangle (in screen space) is visible / not clipped. to perform coarse clipping on user's side.
@[c:'ImGui_GetTime']
fn get_time() f64

// get global imgui time. incremented by io.DeltaTime every frame.
@[c:'ImGui_GetFrameCount']
fn get_frame_count() int

// get global imgui frame count. incremented by 1 every frame.
@[c:'ImGui_GetDrawListSharedData']
fn get_draw_list_shared_data() &C.ImDrawListSharedData

// you may use this when creating your own ImDrawList instances.
@[c:'ImGui_GetStyleColorName']
fn get_style_color_name(idx Col) &i8

// get a string corresponding to the enum value (for display, saving, etc.).
@[c:'ImGui_SetStateStorage']
fn set_state_storage(storage &ImGuiStorage)

// replace current window storage with our own (if you want to manipulate it yourself, typically clear subsection of it)
@[c:'ImGui_GetStateStorage']
fn get_state_storage() &ImGuiStorage

// Text Utilities
@[c:'ImGui_CalcTextSize']
fn calc_text_size(text &i8) ImVec2

// Implied text_end = NULL, hide_text_after_double_hash = false, wrap_width = -1.0f
@[c:'ImGui_CalcTextSizeEx']
fn calc_text_size_ex(text &i8, text_end &i8, hide_text_after_double_hash bool, wrap_width f32) ImVec2

// Color Utilities
@[c:'ImGui_ColorConvertU32ToFloat4']
fn color_convert_u32_to_float4(in_ ImU32) C.ImVec4

@[c:'ImGui_ColorConvertFloat4ToU32']
fn color_convert_float4_to_u32(in_ C.ImVec4) ImU32

@[c:'ImGui_ColorConvertRGBtoHSV']
fn color_convert_rgb_to_hsv(r f32, g f32, b f32, out_h &f32, out_s &f32, out_v &f32)

@[c:'ImGui_ColorConvertHSVtoRGB']
fn color_convert_hsv_to_rgb(h f32, s f32, v f32, out_r &f32, out_g &f32, out_b &f32)

// Inputs Utilities: Keyboard/Mouse/Gamepad
// - the Key enum contains all possible keyboard, mouse and gamepad inputs (e.g. Key_A, Key_MouseLeft, Key_GamepadDpadUp...).
// - (legacy: before v1.87, we used Key to carry native/user indices as defined by each backends. This was obsoleted in 1.87 (2022-02) and completely removed in 1.91.5 (2024-11). See https://github.com/ocornut/imgui/issues/4921)
// - (legacy: any use of Key will assert when key < 512 to detect passing legacy native/user indices)
@[c:'ImGui_IsKeyDown']
fn is_key_down(key Key) bool

// is key being held.
@[c:'ImGui_IsKeyPressed']
fn is_key_pressed(key Key) bool

// Implied repeat = true
@[c:'ImGui_IsKeyPressedEx']
fn is_key_pressed_ex(key Key, repeat bool) bool

// was key pressed (went from !Down to Down)? if repeat=true, uses io.KeyRepeatDelay / KeyRepeatRate
@[c:'ImGui_IsKeyReleased']
fn is_key_released(key Key) bool

// was key released (went from Down to !Down)?
@[c:'ImGui_IsKeyChordPressed']
fn is_key_chord_pressed(key_chord KeyChord) bool

// was key chord (mods + key) pressed, e.g. you can pass 'ImGuiMod_Ctrl | Key_S' as a key-chord. This doesn't do any routing or focus check, please consider using Shortcut() function instead.
@[c:'ImGui_GetKeyPressedAmount']
fn get_key_pressed_amount(key Key, repeat_delay f32, rate f32) int

// uses provided repeat rate/delay. return a count, most often 0 or 1 but might be >1 if RepeatRate is small enough that DeltaTime > RepeatRate
@[c:'ImGui_GetKeyName']
fn get_key_name(key Key) &i8

// [DEBUG] returns English name of the key. Those names are provided for debugging purpose and are not meant to be saved persistently nor compared.
@[c:'ImGui_SetNextFrameWantCaptureKeyboard']
fn set_next_frame_want_capture_keyboard(want_capture_keyboard bool)

// Override io.WantCaptureKeyboard flag next frame (said flag is left for your application to handle, typically when true it instructs your app to ignore inputs). e.g. force capture keyboard when your widget is being hovered. This is equivalent to setting "io.WantCaptureKeyboard = want_capture_keyboard"; after the next NewFrame() call.
// Inputs Utilities: Shortcut Testing & Routing [BETA]
// - KeyChord = a Key + optional Mod_Alt/ImGuiMod_Ctrl/ImGuiMod_Shift/ImGuiMod_Super.
//       Key_C                          // Accepted by functions taking Key or KeyChord arguments)
//       Mod_Ctrl | Key_C          // Accepted by functions taking KeyChord arguments)
//   only Mod_XXX values are legal to combine with an Key. You CANNOT combine two Key values.
// - The general idea is that several callers may register interest in a shortcut, and only one owner gets it.
//      Parent   -> call Shortcut(Ctrl+S)    // When Parent is focused, Parent gets the shortcut.
//        Child1 -> call Shortcut(Ctrl+S)    // When Child1 is focused, Child1 gets the shortcut (Child1 overrides Parent shortcuts)
//        Child2 -> no call                  // When Child2 is focused, Parent gets the shortcut.
//   The whole system is order independent, so if Child1 makes its calls before Parent, results will be identical.
//   This is an important property as it facilitate working with foreign code or larger codebase.
// - To understand the difference:
//   - IsKeyChordPressed() compares mods and call IsKeyPressed() -> function has no side-effect.
//   - Shortcut() submits a route, routes are resolved, if it currently can be routed it calls IsKeyChordPressed() -> function has (desirable) side-effects as it can prevents another call from getting the route.
// - Visualize registered routes in 'Metrics/Debugger->Inputs'.
@[c:'ImGui_Shortcut']
fn shortcut(key_chord KeyChord, flags InputFlags) bool

@[c:'ImGui_SetNextItemShortcut']
fn set_next_item_shortcut(key_chord KeyChord, flags InputFlags)

// Inputs Utilities: Key/Input Ownership [BETA]
// - One common use case would be to allow your items to disable standard inputs behaviors such
//   as Tab or Alt key handling, Mouse Wheel scrolling, etc.
//   e.g. Button(...); SetItemKeyOwner Key_MouseWheelY); to make hovering/activating a button disable wheel for scrolling.
// - Reminder Key enum include access to mouse buttons and gamepad, so key ownership can apply to them.
// - Many related features are still in imgui_internal.h. For instance, most IsKeyXXX()/IsMouseXXX() functions have an owner-id-aware version.
@[c:'ImGui_SetItemKeyOwner']
fn set_item_key_owner(key Key)

// Set key owner to last item ID if it is hovered or active. Equivalent to 'if (IsItemHovered() || IsItemActive()) { SetKeyOwner(key, GetItemID());'.
// Inputs Utilities: Mouse
// - To refer to a mouse button, you may use named enums in your code e.g. MouseButton_Left, MouseButton_Right.
// - You can also use regular integer: it is forever guaranteed that 0=Left, 1=Right, 2=Middle.
// - Dragging operations are only reported after mouse has moved a certain distance away from the initial clicking position (see 'lock_threshold' and 'io.MouseDraggingThreshold')
@[c:'ImGui_IsMouseDown']
fn is_mouse_down(button MouseButton) bool

// is mouse button held?
@[c:'ImGui_IsMouseClicked']
fn is_mouse_clicked(button MouseButton) bool

// Implied repeat = false
@[c:'ImGui_IsMouseClickedEx']
fn is_mouse_clicked_ex(button MouseButton, repeat bool) bool

// did mouse button clicked? (went from !Down to Down). Same as GetMouseClickedCount() == 1.
@[c:'ImGui_IsMouseReleased']
fn is_mouse_released(button MouseButton) bool

// did mouse button released? (went from Down to !Down)
@[c:'ImGui_IsMouseDoubleClicked']
fn is_mouse_double_clicked(button MouseButton) bool

// did mouse button double-clicked? Same as GetMouseClickedCount() == 2. (note that a double-click will also report IsMouseClicked() == true)
@[c:'ImGui_IsMouseReleasedWithDelay']
fn is_mouse_released_with_delay(button MouseButton, delay f32) bool

// delayed mouse release (use very sparingly!). Generally used with 'delay >= io.MouseDoubleClickTime' + combined with a 'io.MouseClickedLastCount==1' test. This is a very rarely used UI idiom, but some apps use this: e.g. MS Explorer single click on an icon to rename.
@[c:'ImGui_GetMouseClickedCount']
fn get_mouse_clicked_count(button MouseButton) int

// return the number of successive mouse-clicks at the time where a click happen (otherwise 0).
@[c:'ImGui_IsMouseHoveringRect']
fn is_mouse_hovering_rect(r_min ImVec2, r_max ImVec2) bool

// Implied clip = true
@[c:'ImGui_IsMouseHoveringRectEx']
fn is_mouse_hovering_rect_ex(r_min ImVec2, r_max ImVec2, clip bool) bool

// is mouse hovering given bounding rect (in screen space). clipped by current clipping settings, but disregarding of other consideration of focus/window ordering/popup-block.
@[c:'ImGui_IsMousePosValid']
fn is_mouse_pos_valid(mouse_pos &ImVec2) bool

// by convention we use (-FLT_MAX,-FLT_MAX) to denote that there is no mouse available
@[c:'ImGui_IsAnyMouseDown']
fn is_any_mouse_down() bool

// [WILL OBSOLETE] is any mouse button held? This was designed for backends, but prefer having backend maintain a mask of held mouse buttons, because upcoming input queue system will make this invalid.
@[c:'ImGui_GetMousePos']
fn get_mouse_pos() ImVec2

// shortcut to ImGui::GetIO().MousePos provided by user, to be consistent with other calls
@[c:'ImGui_GetMousePosOnOpeningCurrentPopup']
fn get_mouse_pos_on_opening_current_popup() ImVec2

// retrieve mouse position at the time of opening popup we have BeginPopup() into (helper to avoid user backing that value themselves)
@[c:'ImGui_IsMouseDragging']
fn is_mouse_dragging(button MouseButton, lock_threshold f32) bool

// is mouse dragging? (uses io.MouseDraggingThreshold if lock_threshold < 0.0f)
@[c:'ImGui_GetMouseDragDelta']
fn get_mouse_drag_delta(button MouseButton, lock_threshold f32) ImVec2

// return the delta from the initial clicking position while the mouse button is pressed or was just released. This is locked and return 0.0f until the mouse moves past a distance threshold at least once (uses io.MouseDraggingThreshold if lock_threshold < 0.0f)
@[c:'ImGui_ResetMouseDragDelta']
fn reset_mouse_drag_delta()

// Implied button = 0
@[c:'ImGui_ResetMouseDragDeltaEx']
fn reset_mouse_drag_delta_ex(button MouseButton)

//
@[c:'ImGui_GetMouseCursor']
fn get_mouse_cursor() MouseCursor

// get desired mouse cursor shape. Important: reset in ImGui::NewFrame(), this is updated during the frame. valid before Render(). If you use software rendering by setting io.MouseDrawCursor ImGui will render those for you
@[c:'ImGui_SetMouseCursor']
fn set_mouse_cursor(cursor_type MouseCursor)

// set desired mouse cursor shape
@[c:'ImGui_SetNextFrameWantCaptureMouse']
fn set_next_frame_want_capture_mouse(want_capture_mouse bool)

// Override io.WantCaptureMouse flag next frame (said flag is left for your application to handle, typical when true it instucts your app to ignore inputs). This is equivalent to setting "io.WantCaptureMouse = want_capture_mouse;" after the next NewFrame() call.
// Clipboard Utilities
// - Also see the LogToClipboard() function to capture GUI into clipboard, or easily output text data to the clipboard.
@[c:'ImGui_GetClipboardText']
fn get_clipboard_text() &i8

@[c:'ImGui_SetClipboardText']
fn set_clipboard_text(text &i8)

// Settings/.Ini Utilities
// - The disk functions are automatically called if io.IniFilename != NULL (default is "imgui.ini").
// - Set io.IniFilename to NULL to load/save manually. Read io.WantSaveIniSettings description about handling .ini saving manually.
// - Important: default value "imgui.ini" is relative to current working dir! Most apps will want to lock this to an absolute path (e.g. same path as executables).
@[c:'ImGui_LoadIniSettingsFromDisk']
fn load_ini_settings_from_disk(ini_filename &i8)

// call after CreateContext() and before the first call to NewFrame(). NewFrame() automatically calls LoadIniSettingsFromDisk(io.IniFilename).
@[c:'ImGui_LoadIniSettingsFromMemory']
fn load_ini_settings_from_memory(ini_data &i8, ini_size usize)

// call after CreateContext() and before the first call to NewFrame() to provide .ini data from your own data source.
@[c:'ImGui_SaveIniSettingsToDisk']
fn save_ini_settings_to_disk(ini_filename &i8)

// this is automatically called (if io.IniFilename is not empty) a few seconds after any modification that should be reflected in the .ini file (and also by DestroyContext).
@[c:'ImGui_SaveIniSettingsToMemory']
fn save_ini_settings_to_memory(out_ini_size &usize) &i8

// return a zero-terminated string with the .ini data which you can save by your own mean. call when io.WantSaveIniSettings is set, then save data by your own mean and clear io.WantSaveIniSettings.
// Debug Utilities
// - Your main debugging friend is the ShowMetricsWindow() function, which is also accessible from Demo->Tools->Metrics Debugger
@[c:'ImGui_DebugTextEncoding']
fn debug_text_encoding(text &i8)

@[c:'ImGui_DebugFlashStyleColor']
fn debug_flash_style_color(idx Col)

@[c:'ImGui_DebugStartItemPicker']
fn debug_start_item_picker()

@[c:'ImGui_DebugCheckVersionAndDataLayout']
fn debug_check_version_and_data_layout(version_str &i8, sz_io usize, sz_style usize, sz_vec2 usize, sz_vec4 usize, sz_drawvert usize, sz_drawidx usize) bool

// This is called by IMGUI_CHECKVERSION() macro.
@[c2v_variadic]
@[c:'ImGui_DebugLog']
fn debug_log(fmt &i8)

// Call via IMGUI_DEBUG_LOG() for maximum stripping in caller code!
@[c:'ImGui_DebugLogV']
fn debug_log_v(fmt &i8, args C.va_list)

// #ifndef IMGUI_DISABLE_DEBUG_TOOLS
// Memory Allocators
// - Those functions are not reliant on the current context.
// - DLL users: heaps and globals are not shared across DLL boundaries! You will need to call SetCurrentContext() + SetAllocatorFunctions()
//   for each static/DLL boundary you are calling from. Read "Context and Memory Allocators" section of imgui.cpp for more details.
@[c:'ImGui_SetAllocatorFunctions']
fn set_allocator_functions(alloc_func MemAllocFunc, free_func MemFreeFunc, user_data voidptr)

@[c:'ImGui_GetAllocatorFunctions']
fn get_allocator_functions(p_alloc_func  MemAllocFunc, p_free_func  MemFreeFunc, p_user_data &voidptr)

@[c:'ImGui_MemAlloc']
fn mem_alloc(size usize) voidptr

@[c:'ImGui_MemFree']
fn mem_free(ptr voidptr)

//-----------------------------------------------------------------------------
// [SECTION] Flags & Enumerations
//-----------------------------------------------------------------------------
// Flags for ImGui::Begin()
// (Those are per-window flags. There are shared flags in ImGuiIO: io.ConfigWindowsResizeFromEdges and io.ConfigWindowsMoveFromTitleBarOnly)
enum WindowFlags_ {
 none = 0
 no_title_bar = 1 << 0
// Disable title-bar
 no_resize = 1 << 1
// Disable user resizing with the lower-right grip
 no_move = 1 << 2
// Disable user moving the window
 no_scrollbar = 1 << 3
// Disable scrollbars (window can still scroll with mouse or programmatically)
 no_scroll_with_mouse = 1 << 4
// Disable user vertically scrolling with mouse wheel. On child window, mouse wheel will be forwarded to the parent unless NoScrollbar is also set.
 no_collapse = 1 << 5
// Disable user collapsing window by double-clicking on it. Also referred to as Window Menu Button (e.g. within a docking node).
 always_auto_resize = 1 << 6
// Resize every window to its content every frame
 no_background = 1 << 7
// Disable drawing background color (WindowBg, etc.) and outside border. Similar as using SetNextWindowBgAlpha(0.0f).
 no_saved_settings = 1 << 8
// Never load/save settings in .ini file
 no_mouse_inputs = 1 << 9
// Disable catching mouse, hovering test with pass through.
 menu_bar = 1 << 10
// Has a menu-bar
 horizontal_scrollbar = 1 << 11
// Allow horizontal scrollbar to appear (off by default). You may use SetNextWindowContentSize(ImVec2(width,0.0f)); prior to calling Begin() to specify width. Read code in imgui_demo in the "Horizontal Scrolling" section.
 no_focus_on_appearing = 1 << 12
// Disable taking focus when transitioning from hidden to visible state
 no_bring_to_front_on_focus = 1 << 13
// Disable bringing window to front when taking focus (e.g. clicking on it or programmatically giving it focus)
 always_vertical_scrollbar = 1 << 14
// Always show vertical scrollbar (even if ContentSize.y < Size.y)
 always_horizontal_scrollbar = 1 << 15
// Always show horizontal scrollbar (even if ContentSize.x < Size.x)
 no_nav_inputs = 1 << 16
// No keyboard/gamepad navigation within the window
 no_nav_focus = 1 << 17
// No focusing toward this window with keyboard/gamepad navigation (e.g. skipped by CTRL+TAB)
 unsaved_document = 1 << 18
// Display a dot next to the title. When used in a tab/docking context, tab is selected when clicking the X + closure is not assumed (will wait for user to stop submitting the tab). Otherwise closure is assumed when pressing the X, so if you keep submitting the tab may reappear at end of tab bar.
 no_nav = 1 << 16 | 1 << 17
 no_decoration = 1 << 0 | 1 << 1 | 1 << 3 | 1 << 5
 no_inputs = 1 << 9 | 1 << 16 | 1 << 17
// [Internal]
 child_window = 1 << 24
// Don't use! For internal use by BeginChild()
 tooltip = 1 << 25
// Don't use! For internal use by BeginTooltip()
 popup = 1 << 26
// Don't use! For internal use by BeginPopup()
 modal = 1 << 27
// Don't use! For internal use by BeginPopupModal()
 child_menu = 1 << 28
// Don't use! For internal use by BeginMenu()
// Obsolete names
 nav_flattened = 1 << 29
// Obsoleted in 1.90.9: Use ChildFlags_NavFlattened in BeginChild() call.
 always_use_window_padding = 1 << 30
// Obsoleted in 1.90.0: Use ChildFlags_AlwaysUseWindowPadding in BeginChild() call.
	
}

// Flags for ImGui::BeginChild()
// (Legacy: bit 0 must always correspond to ChildFlags_Borders to be backward compatible with old API using 'bool border = false'.
// About using AutoResizeX/AutoResizeY flags:
// - May be combined with SetNextWindowSizeConstraints() to set a min/max size for each axis (see "Demo->Child->Auto-resize with Constraints").
// - Size measurement for a given axis is only performed when the child window is within visible boundaries, or is just appearing.
//   - This allows BeginChild() to return false when not within boundaries (e.g. when scrolling), which is more optimal. BUT it won't update its auto-size while clipped.
//     While not perfect, it is a better default behavior as the always-on performance gain is more valuable than the occasional "resizing after becoming visible again" glitch.
//   - You may also use ChildFlags_AlwaysAutoResize to force an update even when child window is not in view.
//     HOWEVER PLEASE UNDERSTAND THAT DOING SO WILL PREVENT BeginChild() FROM EVER RETURNING FALSE, disabling benefits of coarse clipping.
enum ChildFlags_ {
 none = 0
 borders = 1 << 0
// Show an outer border and enable WindowPadding. (IMPORTANT: this is always == 1 == true for legacy reason)
 always_use_window_padding = 1 << 1
// Pad with style.WindowPadding even if no border are drawn (no padding by default for non-bordered child windows because it makes more sense)
 resize_x = 1 << 2
// Allow resize from right border (layout direction). Enable .ini saving (unless WindowFlags_NoSavedSettings passed to window flags)
 resize_y = 1 << 3
// Allow resize from bottom border (layout direction). "
 auto_resize_x = 1 << 4
// Enable auto-resizing width. Read "IMPORTANT: Size measurement" details above.
 auto_resize_y = 1 << 5
// Enable auto-resizing height. Read "IMPORTANT: Size measurement" details above.
 always_auto_resize = 1 << 6
// Combined with AutoResizeX/AutoResizeY. Always measure size even when child is hidden, always return true, always disable clipping optimization! NOT RECOMMENDED.
 frame_style = 1 << 7
// Style the child window like a framed item: use FrameBg, FrameRounding, FrameBorderSize, FramePadding instead of ChildBg, ChildRounding, ChildBorderSize, WindowPadding.
 nav_flattened = 1 << 8
// [BETA] Share focus scope, allow keyboard/gamepad navigation to cross over parent border to this child or between sibling child windows.
// Obsolete names
 border = 1 << 0
// Renamed in 1.91.1 (August 2024) for consistency.
	
}

// Flags for ImGui::PushItemFlag()
// (Those are shared by all items)
enum ItemFlags_ {
 none = 0
// (Default)
 no_tab_stop = 1 << 0
// false    // Disable keyboard tabbing. This is a "lighter" version of ItemFlags_NoNav.
 no_nav = 1 << 1
// false    // Disable any form of focusing (keyboard/gamepad directional navigation and SetKeyboardFocusHere() calls).
 no_nav_default_focus = 1 << 2
// false    // Disable item being a candidate for default focus (e.g. used by title bar items).
 button_repeat = 1 << 3
// false    // Any button-like behavior will have repeat mode enabled (based on io.KeyRepeatDelay and io.KeyRepeatRate values). Note that you can also call IsItemActive() after any button to tell if it is being held.
 auto_close_popups = 1 << 4
// true     // MenuItem()/Selectable() automatically close their parent popup window.
 allow_duplicate_id = 1 << 5
}

// Flags for ImGui::InputText()
// (Those are per-item flags. There are shared flags in ImGuiIO: io.ConfigInputTextCursorBlink and io.ConfigInputTextEnterKeepActive)
enum InputTextFlags_ {
// Basic filters (also see InputTextFlags_CallbackCharFilter)
 none = 0
 chars_decimal = 1 << 0
// Allow 0123456789.+-*/
 chars_hexadecimal = 1 << 1
// Allow 0123456789ABCDEFabcdef
 chars_scientific = 1 << 2
// Allow 0123456789.+-*/eE (Scientific notation input)
 chars_uppercase = 1 << 3
// Turn a..z into A..Z
 chars_no_blank = 1 << 4
// Filter out spaces, tabs
// Inputs
 allow_tab_input = 1 << 5
// Pressing TAB input a '\t' character into the text field
 enter_returns_true = 1 << 6
// Return 'true' when Enter is pressed (as opposed to every time the value was modified). Consider using IsItemDeactivatedAfterEdit() instead!
 escape_clears_all = 1 << 7
// Escape key clears content if not empty, and deactivate otherwise (contrast to default behavior of Escape to revert)
 ctrl_enter_for_new_line = 1 << 8
// In multi-line mode, validate with Enter, add new line with Ctrl+Enter (default is opposite: validate with Ctrl+Enter, add line with Enter).
// Other options
 read_only = 1 << 9
// Read-only mode
 password = 1 << 10
// Password mode, display all characters as '*', disable copy
 always_overwrite = 1 << 11
// Overwrite mode
 auto_select_all = 1 << 12
// Select entire text when first taking mouse focus
 parse_empty_ref_val = 1 << 13
// InputFloat(), InputInt(), InputScalar() etc. only: parse empty string as zero value.
 display_empty_ref_val = 1 << 14
// InputFloat(), InputInt(), InputScalar() etc. only: when value is zero, do not display it. Generally used with InputTextFlags_ParseEmptyRefVal.
 no_horizontal_scroll = 1 << 15
// Disable following the cursor horizontally
 no_undo_redo = 1 << 16
// Disable undo/redo. Note that input text owns the text data while active, if you want to provide your own undo/redo stack you need e.g. to call ClearActiveID().
// Elide display / Alignment
 elide_left = 1 << 17
// When text doesn't fit, elide left side to ensure right side stays visible. Useful for path/filenames. Single-line only!
// Callback features
 callback_completion = 1 << 18
// Callback on pressing TAB (for completion handling)
 callback_history = 1 << 19
// Callback on pressing Up/Down arrows (for history handling)
 callback_always = 1 << 20
// Callback on each iteration. User code may query cursor position, modify text buffer.
 callback_char_filter = 1 << 21
// Callback on character inputs to replace or discard them. Modify 'EventChar' to replace or discard, or return 1 in callback to discard.
 callback_resize = 1 << 22
// Callback on buffer capacity changes request (beyond 'buf_size' parameter value), allowing the string to grow. Notify when the string wants to be resized (for string types which hold a cache of their Size). You will be provided a new BufSize in the callback and NEED to honor it. (see misc/cpp/imgui_stdlib.h for an example of using this)
 callback_edit = 1 << 23
// Callback on any edit. Note that InputText() already returns true on edit + you can always use IsItemEdited(). The callback is useful to manipulate the underlying buffer while focus is active.
	
// Obsolete names
	
}

// Flags for ImGui::TreeNodeEx(), ImGui::CollapsingHeader*()
enum TreeNodeFlags_ {
 none = 0
 selected = 1 << 0
// Draw as selected
 framed = 1 << 1
// Draw frame with background (e.g. for CollapsingHeader)
 allow_overlap = 1 << 2
// Hit testing to allow subsequent widgets to overlap this one
 no_tree_push_on_open = 1 << 3
// Don't do a TreePush() when open (e.g. for CollapsingHeader) = no extra indent nor pushing on ID stack
 no_auto_open_on_log = 1 << 4
// Don't automatically and temporarily open node when Logging is active (by default logging will automatically open tree nodes)
 default_open = 1 << 5
// Default node to be open
 open_on_double_click = 1 << 6
// Open on double-click instead of simple click (default for multi-select unless any _OpenOnXXX behavior is set explicitly). Both behaviors may be combined.
 open_on_arrow = 1 << 7
// Open when clicking on the arrow part (default for multi-select unless any _OpenOnXXX behavior is set explicitly). Both behaviors may be combined.
 leaf = 1 << 8
// No collapsing, no arrow (use as a convenience for leaf nodes).
 bullet = 1 << 9
// Display a bullet instead of arrow. IMPORTANT: node can still be marked open/close if you don't set the _Leaf flag!
 frame_padding = 1 << 10
// Use FramePadding (even for an unframed text node) to vertically align text baseline to regular widget height. Equivalent to calling AlignTextToFramePadding() before the node.
 span_avail_width = 1 << 11
// Extend hit box to the right-most edge, even if not framed. This is not the default in order to allow adding other items on the same line without using AllowOverlap mode.
 span_full_width = 1 << 12
// Extend hit box to the left-most and right-most edges (cover the indent area).
 span_label_width = 1 << 13
// Narrow hit box + narrow hovering highlight, will only cover the label text.
 span_all_columns = 1 << 14
// Frame will span all columns of its container table (label will still fit in current column)
 label_span_all_columns = 1 << 15
// Label will span all columns of its container table
//ImGuiTreeNodeFlags_NoScrollOnOpen     = 1 << 16,  // FIXME: TODO: Disable automatic scroll on TreePop() if node got just open and contents is not visible
 nav_left_jumps_back_here = 1 << 17
// (WIP) Nav: left direction may move to this TreeNode() from any of its child (items submitted between TreeNode and TreePop)
 collapsing_header = 1 << 1 | 1 << 3 | 1 << 4
 allow_item_overlap = 1 << 2
// Renamed in 1.89.7
 span_text_width = 1 << 13
// Renamed in 1.90.7
	
}

// Flags for OpenPopup*(), BeginPopupContext*(), IsPopupOpen() functions.
// - To be backward compatible with older API which took an 'int mouse_button = 1' argument instead of 'ImGuiPopupFlags flags',
//   we need to treat small flags values as a mouse button index, so we encode the mouse button in the first few bits of the flags.
//   It is therefore guaranteed to be legal to pass a mouse button index in PopupFlags.
// - For the same reason, we exceptionally default the PopupFlags argument of BeginPopupContextXXX functions to 1 instead of 0.
//   IMPORTANT: because the default parameter is 1 (= PopupFlags_MouseButtonRight), if you rely on the default parameter
//   and want to use another flag, you need to pass in the PopupFlags_MouseButtonRight flag explicitly.
// - Multiple buttons currently cannot be combined/or-ed in those functions (we could allow it later).
enum PopupFlags_ {
 none = 0
 mouse_button_left = 0
// For BeginPopupContext*(): open on Left Mouse release. Guaranteed to always be == 0 (same as MouseButton_Left)
 mouse_button_right = 1
// For BeginPopupContext*(): open on Right Mouse release. Guaranteed to always be == 1 (same as MouseButton_Right)
 mouse_button_middle = 2
// For BeginPopupContext*(): open on Middle Mouse release. Guaranteed to always be == 2 (same as MouseButton_Middle)
 mouse_button_mask_ = 31
 mouse_button_default_ = 1
 no_reopen = 1 << 5
// For OpenPopup*(), BeginPopupContext*(): don't reopen same popup if already open (won't reposition, won't reinitialize navigation)
//ImGuiPopupFlags_NoReopenAlwaysNavInit = 1 << 6,   // For OpenPopup*(), BeginPopupContext*(): focus and initialize navigation even when not reopening.
 no_open_over_existing_popup = 1 << 7
// For OpenPopup*(), BeginPopupContext*(): don't open if there's already a popup at the same level of the popup stack
 no_open_over_items = 1 << 8
// For BeginPopupContextWindow(): don't return true when hovering items, only when hovering empty space
 any_popup_id = 1 << 10
// For IsPopupOpen(): ignore the ID parameter and test for any popup.
 any_popup_level = 1 << 11
// For IsPopupOpen(): search/test at any level of the popup stack (default test in the current level)
 any_popup = 1 << 10 | 1 << 11
}

// Flags for ImGui::Selectable()
enum SelectableFlags_ {
 none = 0
 no_auto_close_popups = 1 << 0
// Clicking this doesn't close parent popup window (overrides ItemFlags_AutoClosePopups)
 span_all_columns = 1 << 1
// Frame will span all columns of its container table (text will still fit in current column)
 allow_double_click = 1 << 2
// Generate press events on double clicks too
 disabled = 1 << 3
// Cannot be selected, display grayed out text
 allow_overlap = 1 << 4
// (WIP) Hit testing to allow subsequent widgets to overlap this one
 highlight = 1 << 5
// Make the item be displayed as if it is hovered
 dont_close_popups = 1 << 0
// Renamed in 1.91.0
 allow_item_overlap = 1 << 4
// Renamed in 1.89.7
	
}

// Flags for ImGui::BeginCombo()
enum ComboFlags_ {
 none = 0
 popup_align_left = 1 << 0
// Align the popup toward the left by default
 height_small = 1 << 1
// Max ~4 items visible. Tip: If you want your combo popup to be a specific size you can use SetNextWindowSizeConstraints() prior to calling BeginCombo()
 height_regular = 1 << 2
// Max ~8 items visible (default)
 height_large = 1 << 3
// Max ~20 items visible
 height_largest = 1 << 4
// As many fitting items as possible
 no_arrow_button = 1 << 5
// Display on the preview box without the square arrow button
 no_preview = 1 << 6
// Display only a square arrow button
 width_fit_preview = 1 << 7
// Width dynamically calculated from preview contents
 height_mask_ = 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4
}

// Flags for ImGui::BeginTabBar()
enum TabBarFlags_ {
 none = 0
 reorderable = 1 << 0
// Allow manually dragging tabs to re-order them + New tabs are appended at the end of list
 auto_select_new_tabs = 1 << 1
// Automatically select new tabs when they appear
 tab_list_popup_button = 1 << 2
// Disable buttons to open the tab list popup
 no_close_with_middle_mouse_button = 1 << 3
// Disable behavior of closing tabs (that are submitted with p_open != NULL) with middle mouse button. You may handle this behavior manually on user's side with if (IsItemHovered() && IsMouseClicked(2)) *p_open = false.
 no_tab_list_scrolling_buttons = 1 << 4
// Disable scrolling buttons (apply when fitting policy is TabBarFlags_FittingPolicyScroll)
 no_tooltip = 1 << 5
// Disable tooltips when hovering a tab
 draw_selected_overline = 1 << 6
// Draw selected overline markers over selected tab
 fitting_policy_resize_down = 1 << 7
// Resize tabs when they don't fit
 fitting_policy_scroll = 1 << 8
// Add scroll buttons when tabs don't fit
 fitting_policy_mask_ = 1 << 7 | 1 << 8
 fitting_policy_default_ = 1 << 7
}

// Flags for ImGui::BeginTabItem()
enum TabItemFlags_ {
 none = 0
 unsaved_document = 1 << 0
// Display a dot next to the title + set TabItemFlags_NoAssumedClosure.
 set_selected = 1 << 1
// Trigger flag to programmatically make the tab selected when calling BeginTabItem()
 no_close_with_middle_mouse_button = 1 << 2
// Disable behavior of closing tabs (that are submitted with p_open != NULL) with middle mouse button. You may handle this behavior manually on user's side with if (IsItemHovered() && IsMouseClicked(2)) *p_open = false.
 no_push_id = 1 << 3
// Don't call PushID()/PopID() on BeginTabItem()/EndTabItem()
 no_tooltip = 1 << 4
// Disable tooltip for the given tab
 no_reorder = 1 << 5
// Disable reordering this tab or having another tab cross over this tab
 leading = 1 << 6
// Enforce the tab position to the left of the tab bar (after the tab list popup button)
 trailing = 1 << 7
// Enforce the tab position to the right of the tab bar (before the scrolling buttons)
 no_assumed_closure = 1 << 8
}

// Flags for ImGui::IsWindowFocused()
enum FocusedFlags_ {
 none = 0
 child_windows = 1 << 0
// Return true if any children of the window is focused
 root_window = 1 << 1
// Test from root window (top most parent of the current hierarchy)
 any_window = 1 << 2
// Return true if any window is focused. Important: If you are trying to tell how to dispatch your low-level inputs, do NOT use this. Use 'io.WantCaptureMouse' instead! Please read the FAQ!
 no_popup_hierarchy = 1 << 3
// Do not consider popup hierarchy (do not treat popup emitter as parent of popup) (when used with _ChildWindows or _RootWindow)
//ImGuiFocusedFlags_DockHierarchy               = 1 << 4,   // Consider docking hierarchy (treat dockspace host as parent of docked window) (when used with _ChildWindows or _RootWindow)
 root_and_child_windows = 1 << 1 | 1 << 0
}

// Flags for ImGui::IsItemHovered(), ImGui::IsWindowHovered()
// Note: if you are trying to check whether your mouse should be dispatched to Dear ImGui or to your app, you should use 'io.WantCaptureMouse' instead! Please read the FAQ!
// Note: windows with the WindowFlags_NoInputs flag are ignored by IsWindowHovered() calls.
enum HoveredFlags_ {
 none = 0
// Return true if directly over the item/window, not obstructed by another window, not obstructed by an active popup or modal blocking inputs under them.
 child_windows = 1 << 0
// IsWindowHovered() only: Return true if any children of the window is hovered
 root_window = 1 << 1
// IsWindowHovered() only: Test from root window (top most parent of the current hierarchy)
 any_window = 1 << 2
// IsWindowHovered() only: Return true if any window is hovered
 no_popup_hierarchy = 1 << 3
// IsWindowHovered() only: Do not consider popup hierarchy (do not treat popup emitter as parent of popup) (when used with _ChildWindows or _RootWindow)
//ImGuiHoveredFlags_DockHierarchy               = 1 << 4,   // IsWindowHovered() only: Consider docking hierarchy (treat dockspace host as parent of docked window) (when used with _ChildWindows or _RootWindow)
 allow_when_blocked_by_popup = 1 << 5
// Return true even if a popup window is normally blocking access to this item/window
//ImGuiHoveredFlags_AllowWhenBlockedByModal     = 1 << 6,   // Return true even if a modal popup window is normally blocking access to this item/window. FIXME-TODO: Unavailable yet.
 allow_when_blocked_by_active_item = 1 << 7
// Return true even if an active item is blocking access to this item/window. Useful for Drag and Drop patterns.
 allow_when_overlapped_by_item = 1 << 8
// IsItemHovered() only: Return true even if the item uses AllowOverlap mode and is overlapped by another hoverable item.
 allow_when_overlapped_by_window = 1 << 9
// IsItemHovered() only: Return true even if the position is obstructed or overlapped by another window.
 allow_when_disabled = 1 << 10
// IsItemHovered() only: Return true even if the item is disabled
 no_nav_override = 1 << 11
// IsItemHovered() only: Disable using keyboard/gamepad navigation state when active, always query mouse
 allow_when_overlapped = 1 << 8 | 1 << 9
 rect_only = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9
 root_and_child_windows = 1 << 1 | 1 << 0
// Tooltips mode
// - typically used in IsItemHovered() + SetTooltip() sequence.
// - this is a shortcut to pull flags from 'style.HoverFlagsForTooltipMouse' or 'style.HoverFlagsForTooltipNav' where you can reconfigure desired behavior.
//   e.g. 'TooltipHoveredFlagsForMouse' defaults to 'ImGuiHoveredFlags_Stationary | HoveredFlags_DelayShort'.
// - for frequently actioned or hovered items providing a tooltip, you want may to use HoveredFlags_ForTooltip (stationary + delay) so the tooltip doesn't show too often.
// - for items which main purpose is to be hovered, or items with low affordance, or in less consistent apps, prefer no delay or shorter delay.
 for_tooltip = 1 << 12
// Shortcut for standard flags when using IsItemHovered() + SetTooltip() sequence.
// (Advanced) Mouse Hovering delays.
// - generally you can use HoveredFlags_ForTooltip to use application-standardized flags.
// - use those if you need specific overrides.
 stationary = 1 << 13
// Require mouse to be stationary for style.HoverStationaryDelay (~0.15 sec) _at least one time_. After this, can move on same item/window. Using the stationary test tends to reduces the need for a long delay.
 delay_none = 1 << 14
// IsItemHovered() only: Return true immediately (default). As this is the default you generally ignore this.
 delay_short = 1 << 15
// IsItemHovered() only: Return true after style.HoverDelayShort elapsed (~0.15 sec) (shared between items) + requires mouse to be stationary for style.HoverStationaryDelay (once per item).
 delay_normal = 1 << 16
// IsItemHovered() only: Return true after style.HoverDelayNormal elapsed (~0.40 sec) (shared between items) + requires mouse to be stationary for style.HoverStationaryDelay (once per item).
 no_shared_delay = 1 << 17
}

// Flags for ImGui::BeginDragDropSource(), ImGui::AcceptDragDropPayload()
enum DragDropFlags_ {
 none = 0
// BeginDragDropSource() flags
 source_no_preview_tooltip = 1 << 0
// Disable preview tooltip. By default, a successful call to BeginDragDropSource opens a tooltip so you can display a preview or description of the source contents. This flag disables this behavior.
 source_no_disable_hover = 1 << 1
// By default, when dragging we clear data so that IsItemHovered() will return false, to avoid subsequent user code submitting tooltips. This flag disables this behavior so you can still call IsItemHovered() on the source item.
 source_no_hold_to_open_others = 1 << 2
// Disable the behavior that allows to open tree nodes and collapsing header by holding over them while dragging a source item.
 source_allow_null_id = 1 << 3
// Allow items such as Text(), Image() that have no unique identifier to be used as drag source, by manufacturing a temporary identifier based on their window-relative position. This is extremely unusual within the dear imgui ecosystem and so we made it explicit.
 source_extern = 1 << 4
// External source (from outside of dear imgui), won't attempt to read current item/window info. Will always return true. Only one Extern source can be active simultaneously.
 payload_auto_expire = 1 << 5
// Automatically expire the payload if the source cease to be submitted (otherwise payloads are persisting while being dragged)
 payload_no_cross_context = 1 << 6
// Hint to specify that the payload may not be copied outside current dear imgui context.
 payload_no_cross_process = 1 << 7
// Hint to specify that the payload may not be copied outside current process.
// AcceptDragDropPayload() flags
 accept_before_delivery = 1 << 10
// AcceptDragDropPayload() will returns true even before the mouse button is released. You can then call IsDelivery() to test if the payload needs to be delivered.
 accept_no_draw_default_rect = 1 << 11
// Do not draw the default highlight rectangle when hovering over target.
 accept_no_preview_tooltip = 1 << 12
// Request hiding the BeginDragDropSource tooltip from the BeginDragDropTarget site.
 accept_peek_only = 1 << 10 | 1 << 11
// For peeking ahead and inspecting the payload before delivery.
 source_auto_expire_payload = 1 << 5
// Renamed in 1.90.9
	
}

// Standard Drag and Drop payload types. You can define you own payload types using short strings. Types starting with '_' are defined by Dear ImGui.
// float[3]: Standard type for colors, without alpha. User code may use this type.
// float[4]: Standard type for colors. User code may use this type.
// A primary data type
enum DataType_ {
 s8
// signed char / char (with sensible compilers)
 u8
// unsigned char
 s16
// short
 u16
// unsigned short
 s32
// int
 u32
// unsigned int
 s64
// long long / __int64
 u64
// unsigned long long / unsigned __int64
 float
// float
 double
// double
 bool
// bool (provided for user convenience, not supported by scalar widgets)
 string
// char* (provided for user convenience, not supported by scalar widgets)
 count
}

// A cardinal direction

const ( // empty enum
// Forward declared enum type Dir
 dir_none = -1
 dir_left = 0
 dir_right = 1
 dir_up = 2
 dir_down = 3
 dir_count = 5
)

// A sorting direction

const ( // empty enum
// Forward declared enum type SortDirection
 sort_direction_none = 0
 sort_direction_ascending = 1
// Ascending = 0->9, A->Z etc.
 sort_direction_descending = 2
// Descending = 9->0, Z->A etc.
)

// A key identifier  Key_XXX or Mod_XXX value): can represent Keyboard, Mouse and Gamepad values.
// All our named keys are >= 512. Keys value 0 to 511 are left unused and were legacy native/opaque key values (< 1.87).
// Support for legacy keys was completely removed in 1.91.5.
// Read details about the 1.87+ transition : https://github.com/ocornut/imgui/issues/4921
// Note that "Keys" related to physical keys and are not the same concept as input "Characters", the later are submitted via io.AddInputCharacter().
// The keyboard key enum values are named after the keys on a standard US keyboard, and on other keyboard types the keys reported may not match the keycaps.

const ( // empty enum
// Forward declared enum type Key
// Keyboard
 key_none = 0
 key_named_key_begin = 512
// First valid key value (other than 0)
 key_tab = 512
// == Key_NamedKey_BEGIN
 key_left_arrow = 3
 key_right_arrow = 4
 key_up_arrow = 5
 key_down_arrow = 6
 key_page_up = 7
 key_page_down = 8
 key_home = 9
 key_end = 10
 key_insert = 11
 key_delete = 12
 key_backspace = 13
 key_space = 14
 key_enter = 15
 key_escape = 16
 key_left_ctrl = 17
 key_left_shift = 18
 key_left_alt = 19
 key_left_super = 20
 key_right_ctrl = 21
 key_right_shift = 22
 key_right_alt = 23
 key_right_super = 24
 key_menu = 25
 key_0 = 26
 key_1 = 27
 key_2 = 28
 key_3 = 29
 key_4 = 30
 key_5 = 31
 key_6 = 32
 key_7 = 33
 key_8 = 34
 key_9 = 35
 key_a = 36
 key_b = 37
 key_c = 38
 key_d = 39
 key_e = 40
 key_f = 41
 key_g = 42
 key_h = 43
 key_i = 44
 key_j = 45
 key_k = 46
 key_l = 47
 key_m = 48
 key_n = 49
 key_o = 50
 key_p = 51
 key_q = 52
 key_r = 53
 key_s = 54
 key_t = 55
 key_u = 56
 key_v = 57
 key_w = 58
 key_x = 59
 key_y = 60
 key_z = 61
 key_f1 = 62
 key_f2 = 63
 key_f3 = 64
 key_f4 = 65
 key_f5 = 66
 key_f6 = 67
 key_f7 = 68
 key_f8 = 69
 key_f9 = 70
 key_f10 = 71
 key_f11 = 72
 key_f12 = 73
 key_f13 = 74
 key_f14 = 75
 key_f15 = 76
 key_f16 = 77
 key_f17 = 78
 key_f18 = 79
 key_f19 = 80
 key_f20 = 81
 key_f21 = 82
 key_f22 = 83
 key_f23 = 84
 key_f24 = 85
 key_apostrophe = 86
// '
 key_comma = 87
// ,
 key_minus = 88
// -
 key_period = 89
// .
 key_slash = 90
// /
 key_semicolon = 91
// ;
 key_equal = 92
// =
 key_left_bracket = 93
// [
 key_backslash = 94
// \ (this text inhibit multiline comment caused by backslash)
 key_right_bracket = 95
// ]
 key_grave_accent = 96
// `
 key_caps_lock = 97
 key_scroll_lock = 98
 key_num_lock = 99
 key_print_screen = 100
 key_pause = 101
 key_keypad0 = 102
 key_keypad1 = 103
 key_keypad2 = 104
 key_keypad3 = 105
 key_keypad4 = 106
 key_keypad5 = 107
 key_keypad6 = 108
 key_keypad7 = 109
 key_keypad8 = 110
 key_keypad9 = 111
 key_keypad_decimal = 112
 key_keypad_divide = 113
 key_keypad_multiply = 114
 key_keypad_subtract = 115
 key_keypad_add = 116
 key_keypad_enter = 117
 key_keypad_equal = 118
 key_app_back = 119
// Available on some keyboard/mouses. Often referred as "Browser Back"
 key_app_forward = 120
 key_oem102 = 121
// Non-US backslash.
// Gamepad (some of those are analog values, 0.0f to 1.0f)                          // NAVIGATION ACTION
// (download controller mapping PNG/PSD at http://dearimgui.com/controls_sheets)
 key_gamepad_start = 122
// Menu (Xbox)      + (Switch)   Start/Options (PS)
 key_gamepad_back = 123
// View (Xbox)      - (Switch)   Share (PS)
 key_gamepad_face_left = 124
// X (Xbox)         Y (Switch)   Square (PS)        // Tap: Toggle Menu. Hold: Windowing mode (Focus/Move/Resize windows)
 key_gamepad_face_right = 125
// B (Xbox)         A (Switch)   Circle (PS)        // Cancel / Close / Exit
 key_gamepad_face_up = 126
// Y (Xbox)         X (Switch)   Triangle (PS)      // Text Input / On-screen Keyboard
 key_gamepad_face_down = 127
// A (Xbox)         B (Switch)   Cross (PS)         // Activate / Open / Toggle / Tweak
 key_gamepad_dpad_left = 128
// D-pad Left                                       // Move / Tweak / Resize Window (in Windowing mode)
 key_gamepad_dpad_right = 129
// D-pad Right                                      // Move / Tweak / Resize Window (in Windowing mode)
 key_gamepad_dpad_up = 130
// D-pad Up                                         // Move / Tweak / Resize Window (in Windowing mode)
 key_gamepad_dpad_down = 131
// D-pad Down                                       // Move / Tweak / Resize Window (in Windowing mode)
 key_gamepad_l1 = 132
// L Bumper (Xbox)  L (Switch)   L1 (PS)            // Tweak Slower / Focus Previous (in Windowing mode)
 key_gamepad_r1 = 133
// R Bumper (Xbox)  R (Switch)   R1 (PS)            // Tweak Faster / Focus Next (in Windowing mode)
 key_gamepad_l2 = 134
// L Trig. (Xbox)   ZL (Switch)  L2 (PS) [Analog]
 key_gamepad_r2 = 135
// R Trig. (Xbox)   ZR (Switch)  R2 (PS) [Analog]
 key_gamepad_l3 = 136
// L Stick (Xbox)   L3 (Switch)  L3 (PS)
 key_gamepad_r3 = 137
// R Stick (Xbox)   R3 (Switch)  R3 (PS)
 key_gamepad_ls_tick_left = 138
// [Analog]                                         // Move Window (in Windowing mode)
 key_gamepad_ls_tick_right = 139
// [Analog]                                         // Move Window (in Windowing mode)
 key_gamepad_ls_tick_up = 140
// [Analog]                                         // Move Window (in Windowing mode)
 key_gamepad_ls_tick_down = 141
// [Analog]                                         // Move Window (in Windowing mode)
 key_gamepad_rs_tick_left = 142
// [Analog]
 key_gamepad_rs_tick_right = 143
// [Analog]
 key_gamepad_rs_tick_up = 144
// [Analog]
 key_gamepad_rs_tick_down = 145
// [Analog]
// Aliases: Mouse Buttons (auto-submitted from AddMouseButtonEvent() calls)
// - This is mirroring the data also written to io.MouseDown[], io.MouseWheel, in a format allowing them to be accessed via standard key API.
 key_mouse_left = 146
 key_mouse_right = 147
 key_mouse_middle = 148
 key_mouse_x1 = 149
 key_mouse_x2 = 150
 key_mouse_wheel_x = 151
 key_mouse_wheel_y = 152
// [Internal] Reserved for mod storage
 key_reserved_for_mod_ctrl = 153
 key_reserved_for_mod_shift = 154
 key_reserved_for_mod_alt = 155
 key_reserved_for_mod_super = 156
 key_named_key_end = 157
// Keyboard Modifiers (explicitly submitted by backend via AddKeyEvent() calls)
// - This is mirroring the data also written to io.KeyCtrl, io.KeyShift, io.KeyAlt, io.KeySuper, in a format allowing
//   them to be accessed via standard key API, allowing calls such as IsKeyPressed(), IsKeyReleased(), querying duration etc.
// - Code polling every key (e.g. an interface to detect a key press for input mapping) might want to ignore those
//   and prefer using the real keys (e.g. Key_LeftCtrl, Key_RightCtrl instead of Mod_Ctrl).
// - In theory the value of keyboard modifiers should be roughly equivalent to a logical or of the equivalent left/right keys.
//   In practice: it's complicated; mods are often provided from different sources. Keyboard layout, IME, sticky keys and
//   backends tend to interfere and break that equivalence. The safer decision is to relay that ambiguity down to the end-user...
// - On macOS, we swap Cmd(Super) and Ctrl keys at the time of the io.AddKeyEvent() call.
 mod_none = 0
 mod_ctrl = 1 << 12
// Ctrl (non-macOS), Cmd (macOS)
 mod_shift = 1 << 13
// Shift
 mod_alt = 1 << 14
// Option/Menu
 mod_super = 1 << 15
// Windows/Super (non-macOS), Ctrl (macOS)
 mod_mask_ = 61440
// 4-bits
// [Internal] If you need to iterate all keys (for e.g. an input mapper) you may use Key_NamedKey_BEGIN. Key_NamedKey_END.
 key_named_key_count = key_named_key_end - key_named_key_begin
//ImGuiKey_KeysData_SIZE        = Key_NamedKey_COUNT,  // Size of KeysData[]: only hold named keys
//ImGuiKey_KeysData_OFFSET      = Key_NamedKey_BEGIN,  // Accesses to io.KeysData[] must use (key - Key_NamedKey_BEGIN) index.
 key_count = key_named_key_end
// Obsoleted in 1.91.5 because it was extremely misleading (since named keys don't start at 0 anymore)
 mod_shortcut = mod_ctrl
// Removed in 1.90.7, you can now simply use Mod_Ctrl
 key_mod_ctrl = mod_ctrl
 key_mod_shift = mod_shift
 key_mod_alt = mod_alt
 key_mod_super = mod_super
// Renamed in 1.89

//ImGuiKey_KeyPadEnter = Key_KeypadEnter,              // Renamed in 1.87

)

// Flags for Shortcut(), SetNextItemShortcut(),
// (and for upcoming extended versions of IsKeyPressed(), IsMouseClicked(), Shortcut(), SetKeyOwner(), SetItemKeyOwner() that are still in imgui_internal.h)
// Don't mistake with InputTextFlags! (which is for ImGui::InputText() function)
enum InputFlags_ {
 none = 0
 repeat = 1 << 0
// Enable repeat. Return true on successive repeats. Default for legacy IsKeyPressed(). NOT Default for legacy IsMouseClicked(). MUST BE == 1.
// Flags for Shortcut(), SetNextItemShortcut()
// - Routing policies: RouteGlobal+OverActive >> RouteActive or RouteFocused (if owner is active item) >> RouteGlobal+OverFocused >> RouteFocused (if in focused window stack) >> RouteGlobal.
// - Default policy is RouteFocused. Can select only 1 policy among all available.
 route_active = 1 << 10
// Route to active item only.
 route_focused = 1 << 11
// Route to windows in the focus stack (DEFAULT). Deep-most focused window takes inputs. Active item takes inputs over deep-most focused window.
 route_global = 1 << 12
// Global route (unless a focused window or active item registered the route).
 route_always = 1 << 13
// Do not register route, poll keys directly.
// - Routing options
 route_over_focused = 1 << 14
// Option: global route: higher priority than focused route (unless active item in focused route).
 route_over_active = 1 << 15
// Option: global route: higher priority than active item. Unlikely you need to use that: will interfere with every active items, e.g. CTRL+A registered by InputText will be overridden by this. May not be fully honored as user/internal code is likely to always assume they can access keys when active.
 route_unless_bg_focused = 1 << 16
// Option: global route: will not be applied if underlying background/void is focused (== no Dear ImGui windows are focused). Useful for overlay applications.
 route_from_root_window = 1 << 17
// Option: route evaluated from the point of view of root window rather than current window.
// Flags for SetNextItemShortcut()
 tooltip = 1 << 18
}

// Configuration flags stored in io.ConfigFlags. Set by user/application.
enum ConfigFlags_ {
 none = 0
 nav_enable_keyboard = 1 << 0
// Master keyboard navigation enable flag. Enable full Tabbing + directional arrows + space/enter to activate.
 nav_enable_gamepad = 1 << 1
// Master gamepad navigation enable flag. Backend also needs to set BackendFlags_HasGamepad.
 no_mouse = 1 << 4
// Instruct dear imgui to disable mouse inputs and interactions.
 no_mouse_cursor_change = 1 << 5
// Instruct backend to not alter mouse cursor shape and visibility. Use if the backend cursor changes are interfering with yours and you don't want to use SetMouseCursor() to change mouse cursor. You may want to honor requests from imgui by reading GetMouseCursor() yourself instead.
 no_keyboard = 1 << 6
// Instruct dear imgui to disable keyboard inputs and interactions. This is done by ignoring keyboard events and clearing existing states.
// User storage (to allow your backend/engine to communicate to code that may be shared between multiple projects. Those flags are NOT used by core Dear ImGui)
 is_srgb = 1 << 20
// Application is SRGB-aware.
 is_touch_screen = 1 << 21
// Application is using a touch screen instead of a mouse.
 nav_enable_set_mouse_pos = 1 << 2
// [moved/renamed in 1.91.4] -> use bool io.ConfigNavMoveSetMousePos
 nav_no_capture_keyboard = 1 << 3
// [moved/renamed in 1.91.4] -> use bool io.ConfigNavCaptureKeyboard
	
}

// Backend capabilities flags stored in io.BackendFlags. Set by imgui_impl_xxx or custom backend.
enum BackendFlags_ {
 none = 0
 has_gamepad = 1 << 0
// Backend Platform supports gamepad and currently has one connected.
 has_mouse_cursors = 1 << 1
// Backend Platform supports honoring GetMouseCursor() value to change the OS cursor shape.
 has_set_mouse_pos = 1 << 2
// Backend Platform supports io.WantSetMousePos requests to reposition the OS mouse position (only used if io.ConfigNavMoveSetMousePos is set).
 renderer_has_vtx_offset = 1 << 3
}

// Enumeration for PushStyleColor() / PopStyleColor()
enum Col_ {
 text
 text_disabled
 window_bg
// Background of normal windows
 child_bg
// Background of child windows
 popup_bg
// Background of popups, menus, tooltips windows
 border
 border_shadow
 frame_bg
// Background of checkbox, radio button, plot, slider, text input
 frame_bg_hovered
 frame_bg_active
 title_bg
// Title bar
 title_bg_active
// Title bar when focused
 title_bg_lapsed
// Title bar when lapsed
 menu_bar_bg
 scrollbar_bg
 scrollbar_grab
 scrollbar_grab_hovered
 scrollbar_grab_active
 check_mark
// Checkbox tick and RadioButton circle
 slider_grab
 slider_grab_active
 button
 button_hovered
 button_active
 header
// Header* ors are used for CollapsingHeader, TreeNode, Selectable, MenuItem
 header_hovered
 header_active
 separator
 separator_hovered
 separator_active
 resize_grip
// Resize grip in lower-right and lower-left corners of windows.
 resize_grip_hovered
 resize_grip_active
 tab_hovered
// Tab background, when hovered
 tab
// Tab background, when tab-bar is focused & tab is unselected
 tab_selected
// Tab background, when tab-bar is focused & tab is selected
 tab_selected_overline
// Tab horizontal overline, when tab-bar is focused & tab is selected
 tab_dimmed
// Tab background, when tab-bar is unfocused & tab is unselected
 tab_dimmed_selected
// Tab background, when tab-bar is unfocused & tab is selected
 tab_dimmed_selected_overline
//..horizontal overline, when tab-bar is unfocused & tab is selected
 plot_lines
 plot_lines_hovered
 plot_histogram
 plot_histogram_hovered
 table_header_bg
// Table header background
 table_border_strong
// Table outer and header borders (prefer using Alpha=1.0 here)
 table_border_light
// Table inner borders (prefer using Alpha=1.0 here)
 table_row_bg
// Table row background (even rows)
 table_row_bg_alt
// Table row background (odd rows)
 text_link
// Hyperlink or
 text_selected_bg
 drag_drop_target
// Rectangle highlighting a drop target
 nav_cursor
// Color of keyboard/gamepad navigation cursor/rectangle, when visible
 nav_windowing_highlight
// Highlight window when using CTRL+TAB
 nav_windowing_dim_bg
// Darken/orize entire screen behind the CTRL+TAB window list, when active
 modal_window_dim_bg
// Darken/orize entire screen behind a modal window, when one is active
 count

	
}

// Enumeration for PushStyleVar() / PopStyleVar() to temporarily modify the ImGuiStyle structure.
// - The enum only refers to fields of ImGuiStyle which makes sense to be pushed/popped inside UI code.
//   During initialization or between frames, feel free to just poke into ImGuiStyle directly.
// - Tip: Use your programming IDE navigation facilities on the names in the _second column_ below to find the actual members and their description.
//   - In Visual Studio: CTRL+comma ("Edit.GoToAll") can follow symbols inside comments, whereas CTRL+F12 ("Edit.GoToImplementation") cannot.
//   - In Visual Studio w/ Visual Assist installed: ALT+G ("VAssistX.GoToImplementation") can also follow symbols inside comments.
//   - In VS Code, CLion, etc.: CTRL+click can follow symbols inside comments.
// - When changing this enum, you need to update the associated internal table GStyleVarInfo[] accordingly. This is where we link enum values to members offset/type.
enum ImGuiStyleVar_ {
// Enum name -------------------------- // Member in ImGuiStyle structure (see ImGuiStyle for descriptions)
 style_var_alpha
// float     Alpha
 style_var_disabled_alpha
// float     DisabledAlpha
 style_var_window_padding
// ImVec2    WindowPadding
 style_var_window_rounding
// float     WindowRounding
 style_var_window_border_size
// float     WindowBorderSize
 style_var_window_min_size
// ImVec2    WindowMinSize
 style_var_window_title_align
// ImVec2    WindowTitleAlign
 style_var_child_rounding
// float     ChildRounding
 style_var_child_border_size
// float     ChildBorderSize
 style_var_popup_rounding
// float     PopupRounding
 style_var_popup_border_size
// float     PopupBorderSize
 style_var_frame_padding
// ImVec2    FramePadding
 style_var_frame_rounding
// float     FrameRounding
 style_var_frame_border_size
// float     FrameBorderSize
 style_var_item_spacing
// ImVec2    ItemSpacing
 style_var_item_inner_spacing
// ImVec2    ItemInnerSpacing
 style_var_indent_spacing
// float     IndentSpacing
 style_var_cell_padding
// ImVec2    CellPadding
 style_var_scrollbar_size
// float     ScrollbarSize
 style_var_scrollbar_rounding
// float     ScrollbarRounding
 style_var_grab_min_size
// float     GrabMinSize
 style_var_grab_rounding
// float     GrabRounding
 style_var_image_border_size
// float     ImageBorderSize
 style_var_tab_rounding
// float     TabRounding
 style_var_tab_border_size
// float     TabBorderSize
 style_var_tab_bar_border_size
// float     TabBarBorderSize
 style_var_tab_bar_overline_size
// float     TabBarOverlineSize
 style_var_table_angled_headers_angle
// float     TableAngledHeadersAngle
 style_var_table_angled_headers_text_align
// ImVec2  TableAngledHeadersTextAlign
 style_var_button_text_align
// ImVec2    ButtonTextAlign
 style_var_selectable_text_align
// ImVec2    SelectableTextAlign
 style_var_separator_text_border_size
// float     SeparatorTextBorderSize
 style_var_separator_text_align
// ImVec2    SeparatorTextAlign
 style_var_separator_text_padding
// ImVec2    SeparatorTextPadding
 style_var_count
}

// Flags for InvisibleButton() [extended in imgui_internal.h]
enum ButtonFlags_ {
 none = 0
 mouse_button_left = 1 << 0
// React on left mouse button (default)
 mouse_button_right = 1 << 1
// React on right mouse button
 mouse_button_middle = 1 << 2
// React on center mouse button
 mouse_button_mask_ = 1 << 0 | 1 << 1 | 1 << 2
// [Internal]
 enable_nav = 1 << 3
}

// Flags for ColorEdit3() / ColorEdit4() / ColorPicker3() / ColorPicker4() / ColorButton()
enum ColorEditFlags_ {
 none = 0
 no_alpha = 1 << 1
//              // ColorEdit, ColorPicker, ColorButton: ignore Alpha component (will only read 3 components from the input pointer).
 no_picker = 1 << 2
//              // ColorEdit: disable picker when clicking on color square.
 no_options = 1 << 3
//              // ColorEdit: disable toggling options menu when right-clicking on inputs/small preview.
 no_small_preview = 1 << 4
//              // ColorEdit, ColorPicker: disable color square preview next to the inputs. (e.g. to show only the inputs)
 no_inputs = 1 << 5
//              // ColorEdit, ColorPicker: disable inputs sliders/text widgets (e.g. to show only the small preview color square).
 no_tooltip = 1 << 6
//              // ColorEdit, ColorPicker, ColorButton: disable tooltip when hovering the preview.
 no_label = 1 << 7
//              // ColorEdit, ColorPicker: disable display of inline text label (the label is still forwarded to the tooltip and picker).
 no_side_preview = 1 << 8
//              // ColorPicker: disable bigger color preview on right side of the picker, use small color square preview instead.
 no_drag_drop = 1 << 9
//              // ColorEdit: disable drag and drop target. ColorButton: disable drag and drop source.
 no_border = 1 << 10
//              // ColorButton: disable border (which is enforced by default)
// Alpha preview
// - Prior to 1.91.8 (2025/01/21): alpha was made opaque in the preview by default using old name ColorEditFlags_AlphaPreview.
// - We now display the preview as transparent by default. You can use ColorEditFlags_AlphaOpaque to use old behavior.
// - The new flags may be combined better and allow finer controls.
 alpha_opaque = 1 << 11
//              // ColorEdit, ColorPicker, ColorButton: disable alpha in the preview,. Contrary to _NoAlpha it may still be edited when calling ColorEdit4()/ColorPicker4(). For ColorButton() this does the same as _NoAlpha.
 alpha_no_bg = 1 << 12
//              // ColorEdit, ColorPicker, ColorButton: disable rendering a checkerboard background behind transparent color.
 alpha_preview_half = 1 << 13
//              // ColorEdit, ColorPicker, ColorButton: display half opaque / half transparent preview.
// User Options (right-click on widget to change some of them).
 alpha_bar = 1 << 16
//              // ColorEdit, ColorPicker: show vertical alpha bar/gradient in picker.
 hdr = 1 << 19
//              // (WIP) ColorEdit: Currently only disable 0.0f..1.0f limits in RGBA edition (note: you probably want to use ColorEditFlags_Float flag as well).
 display_rgb = 1 << 20
// [Display]    // ColorEdit: override _display_ type among RGB/HSV/Hex. ColorPicker: select any combination using one or more of RGB/HSV/Hex.
 display_hsv = 1 << 21
// [Display]    // "
 display_hex = 1 << 22
// [Display]    // "
 uint8 = 1 << 23
// [DataType]   // ColorEdit, ColorPicker, ColorButton: _display_ values formatted as 0..255.
 float = 1 << 24
// [DataType]   // ColorEdit, ColorPicker, ColorButton: _display_ values formatted as 0.0f..1.0f floats instead of 0..255 integers. No round-trip of value via integers.
 picker_hue_bar = 1 << 25
// [Picker]     // ColorPicker: bar for Hue, rectangle for Sat/Value.
 picker_hue_wheel = 1 << 26
// [Picker]     // ColorPicker: wheel for Hue, triangle for Sat/Value.
 input_rgb = 1 << 27
// [Input]      // ColorEdit, ColorPicker: input and output data in RGB format.
 input_hsv = 1 << 28
// [Input]      // ColorEdit, ColorPicker: input and output data in HSV format.
// Defaults Options. You can set application defaults using SetColorEditOptions(). The intent is that you probably don't want to
// override them in most of your calls. Let the user choose via the option menu and/or call SetColorEditOptions() once during startup.
 default_options_ = 1 << 23 | 1 << 20 | 1 << 27 | 1 << 25
// [Internal] Masks
 alpha_mask_ = 1 << 1 | 1 << 11 | 1 << 12 | 1 << 13
 display_mask_ = 1 << 20 | 1 << 21 | 1 << 22
 data_type_mask_ = 1 << 23 | 1 << 24
 picker_mask_ = 1 << 26 | 1 << 25
 input_mask_ = 1 << 27 | 1 << 28
// Obsolete names
 alpha_preview = 0
// [Removed in 1.91.8] This is the default now. Will display a checkerboard unless ColorEditFlags_AlphaNoBg is set.
	
// #ifndef IMGUI_DISABLE_OBSOLETE_FUNCTIONS
	
}

// Flags for DragFloat(), DragInt(), SliderFloat(), SliderInt() etc.
// We use the same sets of flags for DragXXX() and SliderXXX() functions as the features are the same and it makes it easier to swap them.
// (Those are per-item flags. There is shared behavior flag too: ImGuiIO: io.ConfigDragClickToInputText)
enum SliderFlags_ {
 none = 0
 logarithmic = 1 << 5
// Make the widget logarithmic (linear otherwise). Consider using SliderFlags_NoRoundToFormat with this if using a format-string with small amount of digits.
 no_round_to_format = 1 << 6
// Disable rounding underlying value to match precision of the display format string (e.g. %.3f values are rounded to those 3 digits).
 no_input = 1 << 7
// Disable CTRL+Click or Enter key allowing to input text directly into the widget.
 wrap_around = 1 << 8
// Enable wrapping around from max to min and from min to max. Only supported by DragXXX() functions for now.
 clamp_on_input = 1 << 9
// Clamp value to min/max bounds when input manually with CTRL+Click. By default CTRL+Click allows going out of bounds.
 clamp_zero_range = 1 << 10
// Clamp even if min==max==0.0f. Otherwise due to legacy reason DragXXX functions don't clamp with those values. When your clamping limits are dynamic you almost always want to use it.
 no_speed_tweaks = 1 << 11
// Disable keyboard modifiers altering tweak speed. Useful if you want to alter tweak speed yourself based on your own logic.
 always_clamp = 1 << 9 | 1 << 10
 invalid_mask_ = 1879048207
}

// Identify a mouse button.
// Those values are guaranteed to be stable and we frequently use 0/1 directly. Named enums provided for convenience.
enum MouseButton_ {
 left = 0
 right = 1
 middle = 2
 count = 5
}

// Enumeration for GetMouseCursor()
// User code may request backend to display given cursor by calling SetMouseCursor(), which is why we have some cursors that are marked unused here
enum MouseCursor_ {
 none = -1
 arrow = 0
 text_input
// When hovering over InputText, etc.
 resize_all
// (Unused by Dear ImGui functions)
 resize_ns
// When hovering over a horizontal border
 resize_ew
// When hovering over a vertical border or a column
 resize_nesw
// When hovering over the bottom-left corner of a window
 resize_nwse
// When hovering over the bottom-right corner of a window
 hand
// (Unused by Dear ImGui functions. Use for e.g. hyperlinks)
 wait
// When waiting for something to process/load.
 progress
// When waiting for something to process/load, but application is still interactive.
 not_allowed
// When hovering something with disallowed interaction. Usually a crossed circle.
 count
}

// Enumeration for AddMouseSourceEvent() actual source of Mouse Input data.
// Historically we use "Mouse" terminology everywhere to indicate pointer data, e.g. MousePos, IsMousePressed(), io.AddMousePosEvent()
// But that "Mouse" data can come from different source which occasionally may be useful for application to know about.
// You can submit a change of pointer type using io.AddMouseSourceEvent().

const ( // empty enum
// Forward declared enum type MouseSource
 mouse_source_mouse = 0
// Input is coming from an actual mouse.
 mouse_source_touch_screen = 1
// Input is coming from a touch screen (no hovering prior to initial press, less precise initial press aiming, dual-axis wheeling possible).
 mouse_source_pen = 2
// Input is coming from a pressure/magnetic pen (often used in conjunction with high-sampling rates).
 mouse_source_count = 3
)

// Enumeration for ImGui::SetNextWindow***(), SetWindow***(), SetNextItem***() functions
// Represent a condition.
// Important: Treat as a regular enum! Do NOT combine multiple values using binary operators! All the functions above treat 0 as a shortcut to Cond_Always.
enum Cond_ {
 none = 0
// No ition (always set the variable), same as _Always
 always = 1 << 0
// No ition (always set the variable), same as _None
 once = 1 << 1
// Set the variable once per runtime session (only the first call will succeed)
 first_use_ever = 1 << 2
// Set the variable if the object/window has no persistently saved data (no entry in .ini file)
 appearing = 1 << 3
}

//-----------------------------------------------------------------------------
// [SECTION] Tables API flags and structures  TableFlags, TableColumnFlags, TableRowFlags, TableBgTarget, ImGuiTableSortSpecs, ImGuiTableColumnSortSpecs)
//-----------------------------------------------------------------------------
// Flags for ImGui::BeginTable()
// - Important! Sizing policies have complex and subtle side effects, much more so than you would expect.
//   Read comments/demos carefully + experiment with live demos to get acquainted with them.
// - The DEFAULT sizing policies are:
//    - Default to TableFlags_SizingFixedFit    if ScrollX is on, or if host window has WindowFlags_AlwaysAutoResize.
//    - Default to TableFlags_SizingStretchSame if ScrollX is off.
// - When ScrollX is off:
//    - Table defaults to TableFlags_SizingStretchSame -> all Columns defaults to TableColumnFlags_WidthStretch with same weight.
//    - Columns sizing policy allowed: Stretch (default), Fixed/Auto.
//    - Fixed Columns (if any) will generally obtain their requested width (unless the table cannot fit them all).
//    - Stretch Columns will share the remaining width according to their respective weight.
//    - Mixed Fixed/Stretch columns is possible but has various side-effects on resizing behaviors.
//      The typical use of mixing sizing policies is: any number of LEADING Fixed columns, followed by one or two TRAILING Stretch columns.
//      (this is because the visible order of columns have subtle but necessary effects on how they react to manual resizing).
// - When ScrollX is on:
//    - Table defaults to TableFlags_SizingFixedFit -> all Columns defaults to TableColumnFlags_WidthFixed
//    - Columns sizing policy allowed: Fixed/Auto mostly.
//    - Fixed Columns can be enlarged as needed. Table will show a horizontal scrollbar if needed.
//    - When using auto-resizing (non-resizable) fixed columns, querying the content width to use item right-alignment e.g. SetNextItemWidth(-FLT_MIN) doesn't make sense, would create a feedback loop.
//    - Using Stretch columns OFTEN DOES NOT MAKE SENSE if ScrollX is on, UNLESS you have specified a value for 'inner_width' in BeginTable().
//      If you specify a value for 'inner_width' then effectively the scrolling space is known and Stretch or mixed Fixed/Stretch columns become meaningful again.
// - Read on documentation at the top of imgui_tables.cpp for details.
enum TableFlags_ {
// Features
 none = 0
 resizable = 1 << 0
// Enable resizing columns.
 reorderable = 1 << 1
// Enable reordering columns in header row (need calling TableSetupColumn() + TableHeadersRow() to display headers)
 hideable = 1 << 2
// Enable hiding/disabling columns in context menu.
 sortable = 1 << 3
// Enable sorting. Call TableGetSortSpecs() to obtain sort specs. Also see TableFlags_SortMulti and TableFlags_SortTristate.
 no_saved_settings = 1 << 4
// Disable persisting columns order, width and sort settings in the .ini file.
 context_menu_in_body = 1 << 5
// Right-click on columns body/contents will display table context menu. By default it is available in TableHeadersRow().
// Decorations
 row_bg = 1 << 6
// Set each RowBg color with Col_TableRowBg or Col_TableRowBgAlt (equivalent of calling TableSetBgColor with TableBgFlags_RowBg0 on each row manually)
 borders_inner_h = 1 << 7
// Draw horizontal borders between rows.
 borders_outer_h = 1 << 8
// Draw horizontal borders at the top and bottom.
 borders_inner_v = 1 << 9
// Draw vertical borders between columns.
 borders_outer_v = 1 << 10
// Draw vertical borders on the left and right sides.
 borders_h = 1 << 7 | 1 << 8
// Draw horizontal borders.
 borders_v = 1 << 9 | 1 << 10
// Draw vertical borders.
 borders_inner = 1 << 9 | 1 << 7
// Draw inner borders.
 borders_outer = 1 << 10 | 1 << 8
// Draw outer borders.
 borders = 1 << 9 | 1 << 7 | 1 << 10 | 1 << 8
// Draw all borders.
 no_borders_in_body = 1 << 11
// [ALPHA] Disable vertical borders in columns Body (borders will always appear in Headers). -> May move to style
 no_borders_in_body_until_resize = 1 << 12
// [ALPHA] Disable vertical borders in columns Body until hovered for resize (borders will always appear in Headers). -> May move to style
// Sizing Policy (read above for defaults)
 sizing_fixed_fit = 1 << 13
// Columns default to _WidthFixed or _WidthAuto (if resizable or not resizable), matching contents width.
 sizing_fixed_same = 2 << 13
// Columns default to _WidthFixed or _WidthAuto (if resizable or not resizable), matching the maximum contents width of all columns. Implicitly enable TableFlags_NoKeepColumnsVisible.
 sizing_stretch_prop = 3 << 13
// Columns default to _WidthStretch with default weights proportional to each columns contents widths.
 sizing_stretch_same = 4 << 13
// Columns default to _WidthStretch with default weights all equal, unless overridden by TableSetupColumn().
// Sizing Extra Options
 no_host_extend_x = 1 << 16
// Make outer width auto-fit to columns, overriding outer_size.x value. Only available when ScrollX/ScrollY are disabled and Stretch columns are not used.
 no_host_extend_y = 1 << 17
// Make outer height stop exactly at outer_size.y (prevent auto-extending table past the limit). Only available when ScrollX/ScrollY are disabled. Data below the limit will be clipped and not visible.
 no_keep_columns_visible = 1 << 18
// Disable keeping column always minimally visible when ScrollX is off and table gets too small. Not recommended if columns are resizable.
 precise_widths = 1 << 19
// Disable distributing remainder width to stretched columns (width allocation on a 100-wide table with 3 columns: Without this flag: 33,33,34. With this flag: 33,33,33). With larger number of columns, resizing will appear to be less smooth.
// Clipping
 no_clip = 1 << 20
// Disable clipping rectangle for every individual columns (reduce draw command count, items will be able to overflow into other columns). Generally incompatible with TableSetupScrollFreeze().
// Padding
 pad_outer_x = 1 << 21
// Default if BordersOuterV is on. Enable outermost padding. Generally desirable if you have headers.
 no_pad_outer_x = 1 << 22
// Default if BordersOuterV is off. Disable outermost padding.
 no_pad_inner_x = 1 << 23
// Disable inner padding between columns (double inner padding if BordersOuterV is on, single inner padding if BordersOuterV is off).
// Scrolling
 scroll_x = 1 << 24
// Enable horizontal scrolling. Require 'outer_size' parameter of BeginTable() to specify the container size. Changes default sizing policy. Because this creates a child window, ScrollY is currently generally recommended when using ScrollX.
 scroll_y = 1 << 25
// Enable vertical scrolling. Require 'outer_size' parameter of BeginTable() to specify the container size.
// Sorting
 sort_multi = 1 << 26
// Hold shift when clicking headers to sort on multiple column. TableGetSortSpecs() may return specs where (SpecsCount > 1).
 sort_tristate = 1 << 27
// Allow no sorting, disable default sorting. TableGetSortSpecs() may return specs where (SpecsCount == 0).
// Miscellaneous
 highlight_hovered_column = 1 << 28
// Highlight column headers when hovered (may evolve into a fuller highlight)
// [Internal] Combinations and masks
 sizing_mask_ = 1 << 13 | 2 << 13 | 3 << 13 | 4 << 13
}

// Flags for ImGui::TableSetupColumn()
enum TableColumnFlags_ {
// Input configuration flags
 none = 0
 disabled = 1 << 0
// Overriding/master disable flag: hide column, won't show in context menu (unlike calling TableSetColumnEnabled() which manipulates the user accessible state)
 default_hide = 1 << 1
// Default as a hidden/disabled column.
 default_sort = 1 << 2
// Default as a sorting column.
 width_stretch = 1 << 3
// Column will stretch. Preferable with horizontal scrolling disabled (default if table sizing policy is _SizingStretchSame or _SizingStretchProp).
 width_fixed = 1 << 4
// Column will not stretch. Preferable with horizontal scrolling enabled (default if table sizing policy is _SizingFixedFit and table is resizable).
 no_resize = 1 << 5
// Disable manual resizing.
 no_reorder = 1 << 6
// Disable manual reordering this column, this will also prevent other columns from crossing over this column.
 no_hide = 1 << 7
// Disable ability to hide/disable this column.
 no_clip = 1 << 8
// Disable clipping for this column (all NoClip columns will render in a same draw command).
 no_sort = 1 << 9
// Disable ability to sort on this field (even if TableFlags_Sortable is set on the table).
 no_sort_ascending = 1 << 10
// Disable ability to sort in the ascending direction.
 no_sort_descending = 1 << 11
// Disable ability to sort in the descending direction.
 no_header_label = 1 << 12
// TableHeadersRow() will submit an empty label for this column. Convenient for some small columns. Name will still appear in context menu or in angled headers. You may append into this cell by calling TableSetColumnIndex() right after the TableHeadersRow() call.
 no_header_width = 1 << 13
// Disable header text width contribution to automatic column width.
 prefer_sort_ascending = 1 << 14
// Make the initial sort direction Ascending when first sorting on this column (default).
 prefer_sort_descending = 1 << 15
// Make the initial sort direction Descending when first sorting on this column.
 indent_enable = 1 << 16
// Use current Indent value when entering cell (default for column 0).
 indent_disable = 1 << 17
// Ignore current Indent value when entering cell (default for columns > 0). Indentation changes _within_ the cell will still be honored.
 angled_header = 1 << 18
// TableHeadersRow() will submit an angled header row for this column. Note this will add an extra row.
// Output status flags, read-only via TableGetColumnFlags()
 is_enabled = 1 << 24
// Status: is enabled == not hidden by user/api (referred to as "Hide" in _DefaultHide and _NoHide) flags.
 is_visible = 1 << 25
// Status: is visible == is enabled AND not clipped by scrolling.
 is_sorted = 1 << 26
// Status: is currently part of the sort specs
 is_hovered = 1 << 27
// Status: is hovered by mouse
// [Internal] Combinations and masks
 width_mask_ = 1 << 3 | 1 << 4
 indent_mask_ = 1 << 16 | 1 << 17
 status_mask_ = 1 << 24 | 1 << 25 | 1 << 26 | 1 << 27
 no_direct_resize_ = 1 << 30
}

// Flags for ImGui::TableNextRow()
enum TableRowFlags_ {
 none = 0
 headers = 1 << 0
}

// Enum for ImGui::TableSetBgColor()
// Background colors are rendering in 3 layers:
//  - Layer 0: draw with RowBg0 color if set, otherwise draw with ColumnBg0 if set.
//  - Layer 1: draw with RowBg1 color if set, otherwise draw with ColumnBg1 if set.
//  - Layer 2: draw with CellBg color if set.
// The purpose of the two row/columns layers is to let you decide if a background color change should override or blend with the existing color.
// When using TableFlags_RowBg on the table, each row has the RowBg0 color automatically set for odd/even rows.
// If you set the color of RowBg0 target, your color will override the existing RowBg0 color.
// If you set the color of RowBg1 or ColumnBg1 target, your color will blend over the RowBg0 color.
enum TableBgTarget_ {
 none = 0
 row_bg0 = 1
// Set row background color 0 (generally used for background, automatically set when TableFlags_RowBg is used)
 row_bg1 = 2
// Set row background color 1 (generally used for selection marking)
 cell_bg = 3
}

// Sorting specifications for a table (often handling sort specs for a single column, occasionally more)
// Obtained by calling TableGetSortSpecs().
// When 'SpecsDirty == true' you can sort your data. It will be true with sorting specs have changed since last call, or the first time.
// Make sure to set 'SpecsDirty = false' after sorting, else you may wastefully sort your data every frame!
struct ImGuiTableSortSpecs { 
	specs &ImGuiTableColumnSortSpecs
// Pointer to sort spec array.
	specsCount int
// Sort spec count. Most often 1. May be > 1 when TableFlags_SortMulti is enabled. May be == 0 when TableFlags_SortTristate is enabled.
	specsDirty bool
}
// Sorting specification for one column of a table (sizeof == 12 bytes)
struct ImGuiTableColumnSortSpecs { 
	columnUserID ID
// User id of the column (if specified by a TableSetupColumn() call)
	columnIndex ImS16
// Index of the column
	sortOrder ImS16
// Index within parent ImGuiTableSortSpecs (always stored in order starting from 0, tables sorted on a single criteria will always have a 0 here)
	sortDirection SortDirection
}
//-----------------------------------------------------------------------------
// [SECTION] Helpers: Debug log, memory allocations macros, ImVector<>
//-----------------------------------------------------------------------------
// Extra helpers for C applications
@[c:'ImVector_Construct']
fn im_vector_construct(vector voidptr)

// Construct a zero-size ImVector<> (of any type). This is primarily useful when calling ImFontGlyphRangesBuilder_BuildRanges()
@[c:'ImVector_Destruct']
fn im_vector_destruct(vector voidptr)

// Destruct an ImVector<> (of any type). Important: Frees the vector memory but does not call destructors on contained objects (if they have them)
// Build an ImStr from a regular const char* (no data is copied, so you need to make sure the original char* isn't altered as long as you are using the ImStr).
// #if IMGUI_HAS_IMSTR
// #if defined(IMGUI_HAS_IMSTR)
//-----------------------------------------------------------------------------
// Debug Logging into ShowDebugLogWindow(), tty and more.
//-----------------------------------------------------------------------------
// #ifndef IMGUI_DISABLE_DEBUG_TOOLS
//-----------------------------------------------------------------------------
// IM_MALLOC(), IM_FREE(), IM_NEW(), IM_PLACEMENT_NEW(), IM_DELETE()
// We call C++ constructor on own allocated memory via the placement "new(ptr) Type()" syntax.
// Defining a custom placement new() with a custom parameter allows us to bypass including <new> which on some platforms complains when user has disabled exceptions.
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------
// ImVector<>
// Lightweight std::vector<>-like class to avoid dragging dependencies (also, some implementations of STL with debug enabled are absurdly slow, we bypass it so our code runs fast in debug).
//-----------------------------------------------------------------------------
// - You generally do NOT need to care or use this ever. But we need to make it available in imgui.h because some of our public structures are relying on it.
// - We use std-like naming convention here, which is a little unusual for this codebase.
// - Important: clear() frees memory, resize(0) keep the allocated buffer. We use resize(0) a lot to intentionally recycle allocated buffers across frames and amortize our costs.
// - Important: our implementation does NOT call C++ constructors/destructors, we treat everything as raw data! This is intentional but be extra mindful of that,
//   Do NOT use this class as a std::vector replacement in your own code! Many of the structures used by dear imgui can be safely initialized by a zero-memset.
//-----------------------------------------------------------------------------
struct ImVector_ImWchar { 
	size int
	capacity int
	data &C.ImWchar
}
// Instantiation of ImVector<C.ImWchar>
struct ImVector_ImGuiTextFilter_ImGuiTextRange { 
	size int
	capacity int
	data &ImGuiTextFilter_ImGuiTextRange
}
// Instantiation of ImVector<ImGuiTextFilter_ImGuiTextRange>
struct ImVector_char { 
	size int
	capacity int
	data &i8
}
// Instantiation of ImVector<char>
struct ImVector_ImGuiStoragePair { 
	size int
	capacity int
	data &ImGuiStoragePair
}
// Instantiation of ImVector<ImGuiStoragePair>
struct ImVector_ImGuiSelectionRequest { 
	size int
	capacity int
	data &ImGuiSelectionRequest
}
// Instantiation of ImVector<ImGuiSelectionRequest>
struct ImVector_ImDrawCmd { 
	size int
	capacity int
	data &ImDrawCmd
}
// Instantiation of ImVector<ImDrawCmd>
struct ImVector_ImDrawIdx { 
	size int
	capacity int
	data &ImDrawIdx
}
// Instantiation of ImVector<ImDrawIdx>
struct ImVector_ImDrawChannel { 
	size int
	capacity int
	data &ImDrawChannel
}
// Instantiation of ImVector<ImDrawChannel>
struct ImVector_ImDrawVert { 
	size int
	capacity int
	data &ImDrawVert
}
// Instantiation of ImVector<ImDrawVert>
struct ImVector_ImVec2 { 
	size int
	capacity int
	data &ImVec2
}
// Instantiation of ImVector<ImVec2>
struct ImVector_ImVec4 { 
	size int
	capacity int
	data &C.ImVec4
}
// Instantiation of ImVector<C.ImVec4>
struct ImVector_ImTextureID { 
	size int
	capacity int
	data &ImTextureID
}
// Instantiation of ImVector<ImTextureID>
struct ImVector_ImU8 { 
	size int
	capacity int
	data &ImU8
}
// Instantiation of ImVector<ImU8>
struct ImVector_ImDrawListPtr { 
	size int
	capacity int
	data &&ImDrawList
}
// Instantiation of ImVector<ImDrawList*>
struct ImVector_ImU32 { 
	size int
	capacity int
	data &ImU32
}
// Instantiation of ImVector<ImU32>
struct ImVector_ImFontPtr { 
	size int
	capacity int
	data &&ImFont
}
// Instantiation of ImVector<ImFont*>
struct ImVector_ImFontAtlasCustomRect { 
	size int
	capacity int
	data &ImFontAtlasCustomRect
}
// Instantiation of ImVector<ImFontAtlasCustomRect>
struct ImVector_ImFontConfig { 
	size int
	capacity int
	data &ImFontConfig
}
// Instantiation of ImVector<ImFontConfig>
struct ImVector_float { 
	size int
	capacity int
	data &f32
}
// Instantiation of ImVector<float>
struct ImVector_ImU16 { 
	size int
	capacity int
	data &ImU16
}
// Instantiation of ImVector<ImU16>
struct ImVector_ImFontGlyph { 
	size int
	capacity int
	data &ImFontGlyph
}
// Instantiation of ImVector<ImFontGlyph>
//-----------------------------------------------------------------------------
// [SECTION] ImGuiStyle
//-----------------------------------------------------------------------------
// You may modify the ImGui::GetStyle() main instance during initialization and before NewFrame().
// During the frame, use ImGui::PushStyleVar(ImGuiStyleVar_XXXX)/PopStyleVar() to alter the main style values,
// and ImGui::PushStyleColor Col_XXX)/PopStyleColor() for colors.
//-----------------------------------------------------------------------------
struct ImGuiStyle { 
	alpha f32
// Global alpha applies to everything in Dear ImGui.
	disabledAlpha f32
// Additional alpha multiplier applied by BeginDisabled(). Multiply over current value of Alpha.
	windowPadding ImVec2
// Padding within a window.
	windowRounding f32
// Radius of window corners rounding. Set to 0.0f to have rectangular windows. Large values tend to lead to variety of artifacts and are not recommended.
	windowBorderSize f32
// Thickness of border around windows. Generally set to 0.0f or 1.0f. (Other values are not well tested and more CPU/GPU costly).
	windowBorderHoverPadding f32
// Hit-testing extent outside/inside resizing border. Also extend determination of hovered window. Generally meaningfully larger than WindowBorderSize to make it easy to reach borders.
	windowMinSize ImVec2
// Minimum window size. This is a global setting. If you want to constrain individual windows, use SetNextWindowSizeConstraints().
	windowTitleAlign ImVec2
// Alignment for title bar text. Defaults to (0.0f,0.5f) for left-aligned,vertically centered.
	windowMenuButtonPosition Dir
// Side of the collapsing/docking button in the title bar (None/Left/Right). Defaults to Dir_Left.
	childRounding f32
// Radius of child window corners rounding. Set to 0.0f to have rectangular windows.
	childBorderSize f32
// Thickness of border around child windows. Generally set to 0.0f or 1.0f. (Other values are not well tested and more CPU/GPU costly).
	popupRounding f32
// Radius of popup window corners rounding. (Note that tooltip windows use WindowRounding)
	popupBorderSize f32
// Thickness of border around popup/tooltip windows. Generally set to 0.0f or 1.0f. (Other values are not well tested and more CPU/GPU costly).
	framePadding ImVec2
// Padding within a framed rectangle (used by most widgets).
	frameRounding f32
// Radius of frame corners rounding. Set to 0.0f to have rectangular frame (used by most widgets).
	frameBorderSize f32
// Thickness of border around frames. Generally set to 0.0f or 1.0f. (Other values are not well tested and more CPU/GPU costly).
	itemSpacing ImVec2
// Horizontal and vertical spacing between widgets/lines.
	itemInnerSpacing ImVec2
// Horizontal and vertical spacing between within elements of a composed widget (e.g. a slider and its label).
	cellPadding ImVec2
// Padding within a table cell. Cellpadding.x is locked for entire table. CellPadding.y may be altered between different rows.
	touchExtraPadding ImVec2
// Expand reactive bounding box for touch-based system where touch position is not accurate enough. Unfortunately we don't sort widgets so priority on overlap will always be given to the first widget. So don't grow this too much!
	indentSpacing f32
// Horizontal indentation when e.g. entering a tree node. Generally == (FontSize + FramePadding.x*2).
	columnsMinSpacing f32
// Minimum horizontal spacing between two columns. Preferably > (FramePadding.x + 1).
	scrollbarSize f32
// Width of the vertical scrollbar, Height of the horizontal scrollbar.
	scrollbarRounding f32
// Radius of grab corners for scrollbar.
	grabMinSize f32
// Minimum width/height of a grab box for slider/scrollbar.
	grabRounding f32
// Radius of grabs corners rounding. Set to 0.0f to have rectangular slider grabs.
	logSliderDeadzone f32
// The size in pixels of the dead-zone around zero on logarithmic sliders that cross zero.
	imageBorderSize f32
// Thickness of border around Image() calls.
	tabRounding f32
// Radius of upper corners of a tab. Set to 0.0f to have rectangular tabs.
	tabBorderSize f32
// Thickness of border around tabs.
	tabCloseButtonMinWidthSelected f32
// -1: always visible. 0.0f: visible when hovered. >0.0f: visible when hovered if minimum width.
	tabCloseButtonMinWidthUnselected f32
// -1: always visible. 0.0f: visible when hovered. >0.0f: visible when hovered if minimum width. FLT_MAX: never show close button when unselected.
	tabBarBorderSize f32
// Thickness of tab-bar separator, which takes on the tab active color to denote focus.
	tabBarOverlineSize f32
// Thickness of tab-bar overline, which highlights the selected tab-bar.
	tableAngledHeadersAngle f32
// Angle of angled headers (supported values range from -50.0f degrees to +50.0f degrees).
	tableAngledHeadersTextAlign ImVec2
// Alignment of angled headers within the cell
	colorButtonPosition Dir
// Side of the color button in the ColorEdit4 widget (left/right). Defaults to Dir_Right.
	buttonTextAlign ImVec2
// Alignment of button text when button is larger than text. Defaults to (0.5f, 0.5f) (centered).
	selectableTextAlign ImVec2
// Alignment of selectable text. Defaults to (0.0f, 0.0f) (top-left aligned). It's generally important to keep this left-aligned if you want to lay multiple items on a same line.
	separatorTextBorderSize f32
// Thickness of border in SeparatorText()
	separatorTextAlign ImVec2
// Alignment of text within the separator. Defaults to (0.0f, 0.5f) (left aligned, center).
	separatorTextPadding ImVec2
// Horizontal offset of text from each edge of the separator + spacing on other axis. Generally small values. .y is recommended to be == FramePadding.y.
	displayWindowPadding ImVec2
// Apply to regular windows: amount which we enforce to keep visible when moving near edges of your screen.
	displaySafeAreaPadding ImVec2
// Apply to every windows, menus, popups, tooltips: amount where we avoid displaying contents. Adjust if you cannot see the edges of your screen (e.g. on a TV where scaling has not been configured).
	mouseCursorScale f32
// Scale software rendered mouse cursor (when io.MouseDrawCursor is enabled). We apply per-monitor DPI scaling over this scale. May be removed later.
	antiAliasedLines bool
// Enable anti-aliased lines/borders. Disable if you are really tight on CPU/GPU. Latched at the beginning of the frame (copied to ImDrawList).
	antiAliasedLinesUseTex bool
// Enable anti-aliased lines/borders using textures where possible. Require backend to render with bilinear filtering (NOT point/nearest filtering). Latched at the beginning of the frame (copied to ImDrawList).
	antiAliasedFill bool
// Enable anti-aliased edges around filled shapes (rounded rectangles, circles, etc.). Disable if you are really tight on CPU/GPU. Latched at the beginning of the frame (copied to ImDrawList).
	curveTessellationTol f32
// Tessellation tolerance when using PathBezierCurveTo() without a specific number of segments. Decrease for highly tessellated curves (higher quality, more polygons), increase to reduce quality.
	circleTessellationMaxError f32
// Maximum error (in pixels) allowed when using AddCircle()/AddCircleFilled() or drawing rounded corner rectangles with no explicit segment count specified. Decrease for higher quality but more geometry.
// Colors
	colors [56]C.ImVec4
// Behaviors
// (It is possible to modify those fields mid-frame if specific behavior need it, unlike e.g. configuration fields in ImGuiIO)
	hoverStationaryDelay f32
// Delay for IsItemHovered HoveredFlags_Stationary). Time required to consider mouse stationary.
	hoverDelayShort f32
// Delay for IsItemHovered HoveredFlags_DelayShort). Usually used along with HoverStationaryDelay.
	hoverDelayNormal f32
// Delay for IsItemHovered HoveredFlags_DelayNormal). "
	hoverFlagsForTooltipMouse HoveredFlags
// Default flags when using IsItemHovered HoveredFlags_ForTooltip) or BeginItemTooltip()/SetItemTooltip() while using mouse.
	hoverFlagsForTooltipNav HoveredFlags
}
@[c:'ImGuiStyle_ScaleAllSizes']
fn style_scale_all_sizes(self &ImGuiStyle, scale_factor f32)

//-----------------------------------------------------------------------------
// [SECTION] ImGuiIO
//-----------------------------------------------------------------------------
// Communicate most settings and inputs/outputs to Dear ImGui using this structure.
// Access via ImGui::GetIO(). Read 'Programmer guide' section in .cpp file for general usage.
// It is generally expected that:
// - initialization: backends and user code writes to ImGuiIO.
// - main loop: backends writes to ImGuiIO, user code and imgui code reads from ImGuiIO.
//-----------------------------------------------------------------------------
// Also see ImGui::GetPlatformIO() and ImGuiPlatformIO struct for OS/platform related functions: clipboard, IME etc.
//-----------------------------------------------------------------------------
// [Internal] Storage used by IsKeyDown(), IsKeyPressed() etc functions.
// If prior to 1.87 you used io.KeysDownDuration[] (which was marked as internal), you should use GetKeyData(key)->DownDuration and *NOT* io.KeysData[key]->DownDuration.
struct ImGuiKeyData { 
	down bool
// True for if key is down
	downDuration f32
// Duration the key has been down (<0.0f: not pressed, 0.0f: just pressed, >0.0f: time held)
	downDurationPrev f32
// Last frame duration the key has been down
	analogValue f32
}
struct ImGuiIO { 
//------------------------------------------------------------------
// Configuration                            // Default value
//------------------------------------------------------------------
	configFlags ConfigFlags
// = 0              // See ConfigFlags_ enum. Set by user/application. Keyboard/Gamepad navigation options, etc.
	backendFlags BackendFlags
// = 0              // See BackendFlags_ enum. Set by backend (imgui_impl_xxx files or custom backend) to communicate features supported by the backend.
	displaySize ImVec2
// <unset>          // Main display size, in pixels (generally == GetMainViewport()->Size). May change every frame.
	deltaTime f32
// = 1.0f/60.0f     // Time elapsed since last frame, in seconds. May change every frame.
	iniSavingRate f32
// = 5.0f           // Minimum time between saving positions/sizes to .ini file, in seconds.
	iniFilename &i8
// = "imgui.ini"    // Path to .ini file (important: default "imgui.ini" is relative to current working dir!). Set NULL to disable automatic .ini loading/saving or if you want to manually call LoadIniSettingsXXX() / SaveIniSettingsXXX() functions.
	logFilename &i8
// = "imgui_log.txt"// Path to .log file (default parameter to ImGui::LogToFile when no file is specified).
	userData voidptr
// = NULL           // Store your own data.
// Font system
	fonts &ImFontAtlas
// <auto>           // Font atlas: load, rasterize and pack one or more fonts into a single texture.
	fontGlobalScale f32
// = 1.0f           // Global scale all fonts
	fontAllowUserScaling bool
// = false          // [OBSOLETE] Allow user scaling text of individual window with CTRL+Wheel.
	fontDefault &ImFont
// = NULL           // Font to use on NewFrame(). Use NULL to uses Fonts->Fonts[0].
	displayFramebufferScale ImVec2
// = (1, 1)         // For retina display or other situations where window coordinates are different from framebuffer coordinates. This generally ends up in ImDrawData::FramebufferScale.
// Keyboard/Gamepad Navigation options
	configNavSwapGamepadButtons bool
// = false          // Swap Activate<>Cancel (A<>B) buttons, matching typical "Nintendo/Japanese style" gamepad layout.
	configNavMoveSetMousePos bool
// = false          // Directional/tabbing navigation teleports the mouse cursor. May be useful on TV/console systems where moving a virtual mouse is difficult. Will update io.MousePos and set io.WantSetMousePos=true.
	configNavCaptureKeyboard bool
// = true           // Sets io.WantCaptureKeyboard when io.NavActive is set.
	configNavEscapeClearFocusItem bool
// = true           // Pressing Escape can clear focused item + navigation id/highlight. Set to false if you want to always keep highlight on.
	configNavEscapeClearFocusWindow bool
// = false          // Pressing Escape can clear focused window as well (super set of io.ConfigNavEscapeClearFocusItem).
	configNavCursorVisibleAuto bool
// = true           // Using directional navigation key makes the cursor visible. Mouse click hides the cursor.
	configNavCursorVisibleAlways bool
// = false          // Navigation cursor is always visible.
// Miscellaneous options
// (you can visualize and interact with all options in 'Demo->Configuration')
	mouseDrawCursor bool
// = false          // Request ImGui to draw a mouse cursor for you (if you are on a platform without a mouse cursor). Cannot be easily renamed to 'io.ConfigXXX' because this is frequently used by backend implementations.
	configMacOSXBehaviors bool
// = defined(__APPLE__) // Swap Cmd<>Ctrl keys + OS X style text editing cursor movement using Alt instead of Ctrl, Shortcuts using Cmd/Super instead of Ctrl, Line/Text Start and End using Cmd+Arrows instead of Home/End, Double click selects by word instead of selecting whole text, Multi-selection in lists uses Cmd/Super instead of Ctrl.
	configInputTrickleEventQueue bool
// = true           // Enable input queue trickling: some types of events submitted during the same frame (e.g. button down + up) will be spread over multiple frames, improving interactions with low framerates.
	configInputTextCursorBlink bool
// = true           // Enable blinking cursor (optional as some users consider it to be distracting).
	configInputTextEnterKeepActive bool
// = false          // [BETA] Pressing Enter will keep item active and select contents (single-line only).
	configDragClickToInputText bool
// = false          // [BETA] Enable turning DragXXX widgets into text input with a simple mouse click-release (without moving). Not desirable on devices without a keyboard.
	configWindowsResizeFromEdges bool
// = true           // Enable resizing of windows from their edges and from the lower-left corner. This requires BackendFlags_HasMouseCursors for better mouse cursor feedback. (This used to be a per-window WindowFlags_ResizeFromAnySide flag)
	configWindowsMoveFromTitleBarOnly bool
// = false      // Enable allowing to move windows only when clicking on their title bar. Does not apply to windows without a title bar.
	configWindowsCopyContentsWithCtrlC bool
// = false      // [EXPERIMENTAL] CTRL+C copy the contents of focused window into the clipboard. Experimental because: (1) has known issues with nested Begin/End pairs (2) text output quality varies (3) text output is in submission order rather than spatial order.
	configScrollbarScrollByPage bool
// = true           // Enable scrolling page by page when clicking outside the scrollbar grab. When disabled, always scroll to clicked location. When enabled, Shift+Click scrolls to clicked location.
	configMemoryCompactTimer f32
// = 60.0f          // Timer (in seconds) to free transient windows/tables memory buffers when unused. Set to -1.0f to disable.
// Inputs Behaviors
// (other variables, ones which are expected to be tweaked within UI code, are exposed in ImGuiStyle)
	mouseDoubleClickTime f32
// = 0.30f          // Time for a double-click, in seconds.
	mouseDoubleClickMaxDist f32
// = 6.0f           // Distance threshold to stay in to validate a double-click, in pixels.
	mouseDragThreshold f32
// = 6.0f           // Distance threshold before considering we are dragging.
	keyRepeatDelay f32
// = 0.275f         // When holding a key/button, time before it starts repeating, in seconds (for buttons in Repeat mode, etc.).
	keyRepeatRate f32
// = 0.050f         // When holding a key/button, rate at which it repeats, in seconds.
//------------------------------------------------------------------
// Debug options
//------------------------------------------------------------------
// Options to configure Error Handling and how we handle recoverable errors [EXPERIMENTAL]
// - Error recovery is provided as a way to facilitate:
//    - Recovery after a programming error (native code or scripting language - the later tends to facilitate iterating on code while running).
//    - Recovery after running an exception handler or any error processing which may skip code after an error has been detected.
// - Error recovery is not perfect nor guaranteed! It is a feature to ease development.
//   You not are not supposed to rely on it in the course of a normal application run.
// - Functions that support error recovery are using IM_ASSERT_USER_ERROR() instead of IM_ASSERT().
// - By design, we do NOT allow error recovery to be 100% silent. One of the three options needs to be checked!
// - Always ensure that on programmers seats you have at minimum Asserts or Tooltips enabled when making direct imgui API calls!
//   Otherwise it would severely hinder your ability to catch and correct mistakes!
// Read https://github.com/ocornut/imgui/wiki/Error-Handling for details.
// - Programmer seats: keep asserts (default), or disable asserts and keep error tooltips (new and nice!)
// - Non-programmer seats: maybe disable asserts, but make sure errors are resurfaced (tooltips, visible log entries, use callback etc.)
// - Recovery after error/exception: record stack sizes with ErrorRecoveryStoreState(), disable assert, set log callback (to e.g. trigger high-level breakpoint), recover with ErrorRecoveryTryToRecoverState(), restore settings.
	configErrorRecovery bool
// = true       // Enable error recovery support. Some errors won't be detected and lead to direct crashes if recovery is disabled.
	configErrorRecoveryEnableAssert bool
// = true       // Enable asserts on recoverable error. By default call IM_ASSERT() when returning from a failing IM_ASSERT_USER_ERROR()
	configErrorRecoveryEnableDebugLog bool
// = true       // Enable debug log output on recoverable errors.
	configErrorRecoveryEnableTooltip bool
// = true       // Enable tooltip on recoverable errors. The tooltip include a way to enable asserts if they were disabled.
// Option to enable various debug tools showing buttons that will call the IM_DEBUG_BREAK() macro.
// - The Item Picker tool will be available regardless of this being enabled, in order to maximize its discoverability.
// - Requires a debugger being attached, otherwise IM_DEBUG_BREAK() options will appear to crash your application.
//   e.g. io.ConfigDebugIsDebuggerPresent = ::IsDebuggerPresent() on Win32, or refer to ImOsIsDebuggerPresent() imgui_test_engine/imgui_te_utils.cpp for a Unix compatible version).
	configDebugIsDebuggerPresent bool
// = false          // Enable various tools calling IM_DEBUG_BREAK().
// Tools to detect code submitting items with conflicting/duplicate IDs
// - Code should use PushID()/PopID() in loops, or append "##xx" to same-label identifiers.
// - Empty label e.g. Button("") == same ID as parent widget/node. Use Button("##xx") instead!
// - See FAQ https://github.com/ocornut/imgui/blob/master/docs/FAQ.md#q-about-the-id-stack-system
	configDebugHighlightIdConflicts bool
// = true           // Highlight and show an error message popup when multiple items have conflicting identifiers.
	configDebugHighlightIdConflictsShowItemPicker bool
//=true // Show "Item Picker" button in aforementioned popup.
// Tools to test correct Begin/End and BeginChild/EndChild behaviors.
// - Presently Begin()/End() and BeginChild()/EndChild() needs to ALWAYS be called in tandem, regardless of return value of BeginXXX()
// - This is inconsistent with other BeginXXX functions and create confusion for many users.
// - We expect to update the API eventually. In the meanwhile we provide tools to facilitate checking user-code behavior.
	configDebugBeginReturnValueOnce bool
// = false          // First-time calls to Begin()/BeginChild() will return false. NEEDS TO BE SET AT APPLICATION BOOT TIME if you don't want to miss windows.
	configDebugBeginReturnValueLoop bool
// = false          // Some calls to Begin()/BeginChild() will return false. Will cycle through window depths then repeat. Suggested use: add "io.ConfigDebugBeginReturnValue = io.KeyShift" in your main loop then occasionally press SHIFT. Windows should be flickering while running.
// Option to deactivate io.AddFocusEvent(false) handling.
// - May facilitate interactions with a debugger when focus loss leads to clearing inputs data.
// - Backends may have other side-effects on focus loss, so this will reduce side-effects but not necessary remove all of them.
	configDebugIgnoreFocusLoss bool
// = false          // Ignore io.AddFocusEvent(false), consequently not calling io.ClearInputKeys()/io.ClearInputMouse() in input processing.
// Option to audit .ini data
	configDebugIniSettings bool
// = false          // Save .ini data with extra comments (particularly helpful for Docking, but makes saving slower)
//------------------------------------------------------------------
// Platform Identifiers
// (the imgui_impl_xxxx backend files are setting those up for you)
//------------------------------------------------------------------
// Nowadays those would be stored in ImGuiPlatformIO but we are leaving them here for legacy reasons.
// Optional: Platform/Renderer backend name (informational only! will be displayed in About Window) + User data for backend/wrappers to store their own stuff.
	backendPlatformName &i8
// = NULL
	backendRendererName &i8
// = NULL
	backendPlatformUserData voidptr
// = NULL           // User data for platform backend
	backendRendererUserData voidptr
// = NULL           // User data for renderer backend
	backendLanguageUserData voidptr
// = NULL           // User data for non C++ programming language backend
//------------------------------------------------------------------
// Input - Call before calling NewFrame()
//------------------------------------------------------------------
//------------------------------------------------------------------
// Output - Updated by NewFrame() or EndFrame()/Render()
// (when reading from the io.WantCaptureMouse, io.WantCaptureKeyboard flags to dispatch your inputs, it is
//  generally easier and more correct to use their state BEFORE calling NewFrame(). See FAQ for details!)
//------------------------------------------------------------------
	wantCaptureMouse bool
// Set when Dear ImGui will use mouse inputs, in this case do not dispatch them to your main game/application (either way, always pass on mouse inputs to imgui). (e.g. unclicked mouse is hovering over an imgui window, widget is active, mouse was clicked over an imgui window, etc.).
	wantCaptureKeyboard bool
// Set when Dear ImGui will use keyboard inputs, in this case do not dispatch them to your main game/application (either way, always pass keyboard inputs to imgui). (e.g. InputText active, or an imgui window is focused and navigation is enabled, etc.).
	wantTextInput bool
// Mobile/console: when set, you may display an on-screen keyboard. This is set by Dear ImGui when it wants textual keyboard input to happen (e.g. when a InputText widget is active).
	wantSetMousePos bool
// MousePos has been altered, backend should reposition mouse on next frame. Rarely used! Set only when io.ConfigNavMoveSetMousePos is enabled.
	wantSaveIniSettings bool
// When manual .ini load/save is active (io.IniFilename == NULL), this will be set to notify your application that you can call SaveIniSettingsToMemory() and save yourself. Important: clear io.WantSaveIniSettings yourself after saving!
	navActive bool
// Keyboard/Gamepad navigation is currently allowed (will handle Key_NavXXX events) = a window is focused and it doesn't use the WindowFlags_NoNavInputs flag.
	navVisible bool
// Keyboard/Gamepad navigation highlight is visible and allowed (will handle Key_NavXXX events).
	framerate f32
// Estimate of application framerate (rolling average over 60 frames, based on io.DeltaTime), in frame per second. Solely for convenience. Slow applications may not want to use a moving average or may want to reset underlying buffers occasionally.
	metricsRenderVertices int
// Vertices output during last call to Render()
	metricsRenderIndices int
// Indices output during last call to Render() = number of triangles * 3
	metricsRenderWindows int
// Number of visible windows
	metricsActiveWindows int
// Number of active windows
	mouseDelta ImVec2
// Mouse delta. Note that this is zero if either current or previous position are invalid (-FLT_MAX,-FLT_MAX), so a disappearing/reappearing mouse won't have a huge delta.
//------------------------------------------------------------------
// [Internal] Dear ImGui will maintain those fields. Forward compatibility not guaranteed!
//------------------------------------------------------------------
	ctx &C.ImGuiContext
// Parent UI context (needs to be set explicitly by parent).
// Main Input State
// (this block used to be written by backend, since 1.87 it is best to NOT write to those directly, call the AddXXX functions above instead)
// (reading from those variables is fair game, as they are extremely unlikely to be moving anywhere)
	mousePos ImVec2
// Mouse position, in pixels. Set to ImVec2(-FLT_MAX, -FLT_MAX) if mouse is unavailable (on another screen, etc.)
	mouseDown [5]bool
// Mouse buttons: 0=left, 1=right, 2=middle + extras  MouseButton_COUNT == 5). Dear ImGui mostly uses left and right buttons. Other buttons allow us to track if the mouse is being used by your application + available to user as a convenience via IsMouse** API.
	mouseWheel f32
// Mouse wheel Vertical: 1 unit scrolls about 5 lines text. >0 scrolls Up, <0 scrolls Down. Hold SHIFT to turn vertical scroll into horizontal scroll.
	mouseWheelH f32
// Mouse wheel Horizontal. >0 scrolls Left, <0 scrolls Right. Most users don't have a mouse with a horizontal wheel, may not be filled by all backends.
	mouseSource MouseSource
// Mouse actual input peripheral (Mouse/TouchScreen/Pen).
	keyCtrl bool
// Keyboard modifier down: Control
	keyShift bool
// Keyboard modifier down: Shift
	keyAlt bool
// Keyboard modifier down: Alt
	keySuper bool
// Keyboard modifier down: Cmd/Super/Windows
// Other state maintained from data above + IO function calls
	keyMods KeyChord
// Key mods flags (any of Mod_Ctrl/ImGuiMod_Shift/ImGuiMod_Alt/ImGuiMod_Super flags, same as io.KeyCtrl/KeyShift/KeyAlt/KeySuper but merged into flags. Read-only, updated by NewFrame()
	keysData [155]ImGuiKeyData
// Key state for all known keys. Use IsKeyXXX() functions to access this.
	wantCaptureMouseUnlessPopupClose bool
// Alternative to WantCaptureMouse: (WantCaptureMouse == true && WantCaptureMouseUnlessPopupClose == false) when a click over void is expected to close a popup.
	mousePosPrev ImVec2
// Previous mouse position (note that MouseDelta is not necessary == MousePos-MousePosPrev, in case either position is invalid)
	mouseClickedPos [5]ImVec2
// Position at time of clicking
	mouseClickedTime [5]f64
// Time of last click (used to figure out double-click)
	mouseClicked [5]bool
// Mouse button went from !Down to Down (same as MouseClickedCount[x] != 0)
	mouseDoubleClicked [5]bool
// Has mouse button been double-clicked? (same as MouseClickedCount[x] == 2)
	mouseClickedCount [5]ImU16
// == 0 (not clicked), == 1 (same as MouseClicked[]), == 2 (double-clicked), == 3 (triple-clicked) etc. when going from !Down to Down
	mouseClickedLastCount [5]ImU16
// Count successive number of clicks. Stays valid after mouse release. Reset after another click is done.
	mouseReleased [5]bool
// Mouse button went from Down to !Down
	mouseReleasedTime [5]f64
// Time of last released (rarely used! but useful to handle delayed single-click when trying to disambiguate them from double-click).
	mouseDownOwned [5]bool
// Track if button was clicked inside a dear imgui window or over void blocked by a popup. We don't request mouse capture from the application if click started outside ImGui bounds.
	mouseDownOwnedUnlessPopupClose [5]bool
// Track if button was clicked inside a dear imgui window.
	mouseWheelRequestAxisSwap bool
// On a non-Mac system, holding SHIFT requests WheelY to perform the equivalent of a WheelX event. On a Mac system this is already enforced by the system.
	mouseCtrlLeftAsRightClick bool
// (OSX) Set to true when the current click was a Ctrl+click that spawned a simulated right click
	mouseDownDuration [5]f32
// Duration the mouse button has been down (0.0f == just clicked)
	mouseDownDurationPrev [5]f32
// Previous time the mouse button has been down
	mouseDragMaxDistanceSqr [5]f32
// Squared maximum distance of how much mouse has traveled from the clicking point (used for moving thresholds)
	penPressure f32
// Touch/Pen pressure (0.0f to 1.0f, should be >0.0f only when MouseDown[0] == true). Helper storage currently unused by Dear ImGui.
	appFocusLost bool
// Only modify via AddFocusEvent()
	appAcceptingEvents bool
// Only modify via SetAppAcceptingEvents()
	inputQueueSurrogate ImWchar16
// For AddInputCharacterUTF16()
	inputQueueCharacters ImVector_ImWchar
// Queue of _characters_ input (obtained by platform backend). Fill using AddInputCharacter() helper.
// Legacy: before 1.87, we required backend to fill io.KeyMap[] (imgui->native map) during initialization and io.KeysDown[] (native indices) every frame.
// This is still temporarily supported as a legacy feature. However the new preferred scheme is for backend to call io.AddKeyEvent().
//   Old (<1.87):  ImGui::IsKeyPressed(ImGui::GetIO().KeyMap Key_Space]) --> New (1.87+) ImGui::IsKeyPressed Key_Space)
//   Old (<1.87):  ImGui::IsKeyPressed(MYPLATFORM_KEY_SPACE)                  --> New (1.87+) ImGui::IsKeyPressed Key_Space)
// Read https://github.com/ocornut/imgui/issues/4921 for details.
//int       KeyMap Key_COUNT];             // [LEGACY] Input: map of indices into the KeysDown[512] entries array which represent your "native" keyboard state. The first 512 are now unused and should be kept zero. Legacy backend will write into KeyMap[] using Key_ indices which are always >512.
//bool      KeysDown Key_COUNT];           // [LEGACY] Input: Keyboard keys that are pressed (ideally left in the "native" order your engine has access to keyboard keys, so you can use your own defines/enums for keys). This used to be [512] sized. It is now Key_COUNT to allow legacy io.KeysDown[GetKeyIndex(...)] to work without an overflow.
//float     NavInputs NavInput_COUNT];     // [LEGACY] Since 1.88, NavInputs[] was removed. Backends from 1.60 to 1.86 won't build. Feed gamepad inputs via io.AddKeyEvent() and Key_GamepadXXX enums.
//void*     ImeWindowHandle;                    // [Obsoleted in 1.87] Set ImGuiViewport::PlatformHandleRaw instead. Set this to your HWND to get automatic IME cursor positioning.
// Legacy: before 1.91.1, clipboard functions were stored in ImGuiIO instead of ImGuiPlatformIO.
// As this is will affect all users of custom engines/backends, we are providing proper legacy redirection (will obsolete).
	getClipboardTextFn fn (voidptr) &i8
	setClipboardTextFn fn (voidptr, &i8)
	clipboardUserData voidptr
}
// Input Functions
@[c:'ImGuiIO_AddKeyEvent']
fn io_add_key_event(self &ImGuiIO, key Key, down bool)

// Queue a new key down/up event. Key should be "translated" (as in, generally Key_A matches the key end-user would use to emit an 'A' character)
@[c:'ImGuiIO_AddKeyAnalogEvent']
fn io_add_key_analog_event(self &ImGuiIO, key Key, down bool, v f32)

// Queue a new key down/up event for analog values (e.g. Key_Gamepad_ values). Dead-zones should be handled by the backend.
@[c:'ImGuiIO_AddMousePosEvent']
fn io_add_mouse_pos_event(self &ImGuiIO, x f32, y f32)

// Queue a mouse position update. Use -FLT_MAX,-FLT_MAX to signify no mouse (e.g. app not focused and not hovered)
@[c:'ImGuiIO_AddMouseButtonEvent']
fn io_add_mouse_button_event(self &ImGuiIO, button int, down bool)

// Queue a mouse button change
@[c:'ImGuiIO_AddMouseWheelEvent']
fn io_add_mouse_wheel_event(self &ImGuiIO, wheel_x f32, wheel_y f32)

// Queue a mouse wheel update. wheel_y<0: scroll down, wheel_y>0: scroll up, wheel_x<0: scroll right, wheel_x>0: scroll left.
@[c:'ImGuiIO_AddMouseSourceEvent']
fn io_add_mouse_source_event(self &ImGuiIO, source MouseSource)

// Queue a mouse source change (Mouse/TouchScreen/Pen)
@[c:'ImGuiIO_AddFocusEvent']
fn io_add_focus_event(self &ImGuiIO, focused bool)

// Queue a gain/loss of focus for the application (generally based on OS/platform focus of your window)
@[c:'ImGuiIO_AddInputCharacter']
fn io_add_input_character(self &ImGuiIO, c u32)

// Queue a new character input
@[c:'ImGuiIO_AddInputCharacterUTF16']
fn io_add_input_character_utf_16(self &ImGuiIO, c ImWchar16)

// Queue a new character input from a UTF-16 character, it can be a surrogate
@[c:'ImGuiIO_AddInputCharactersUTF8']
fn io_add_input_characters_utf_8(self &ImGuiIO, str &i8)

// Queue a new characters input from a UTF-8 string
@[c:'ImGuiIO_SetKeyEventNativeData']
fn io_set_key_event_native_data(self &ImGuiIO, key Key, native_keycode int, native_scancode int)

// Implied native_legacy_index = -1
@[c:'ImGuiIO_SetKeyEventNativeDataEx']
fn io_set_key_event_native_data_ex(self &ImGuiIO, key Key, native_keycode int, native_scancode int, native_legacy_index int)

// [Optional] Specify index for legacy <1.87 IsKeyXXX() functions with native indices + specify native keycode, scancode.
@[c:'ImGuiIO_SetAppAcceptingEvents']
fn io_set_app_accepting_events(self &ImGuiIO, accepting_events bool)

// Set master flag for accepting key/mouse/text events (default to true). Useful if you have native dialog boxes that are interrupting your application loop/refresh, and you want to disable events being queued while your app is frozen.
@[c:'ImGuiIO_ClearEventsQueue']
fn io_clear_events_queue(self &ImGuiIO)

// Clear all incoming events.
@[c:'ImGuiIO_ClearInputKeys']
fn io_clear_input_keys(self &ImGuiIO)

// Clear current keyboard/gamepad state + current frame text input buffer. Equivalent to releasing all keys/buttons.
@[c:'ImGuiIO_ClearInputMouse']
fn io_clear_input_mouse(self &ImGuiIO)

// Clear current mouse state.
@[c:'ImGuiIO_ClearInputCharacters']
fn io_clear_input_characters(self &ImGuiIO)

// [Obsoleted in 1.89.8] Clear the current frame text input buffer. Now included within ClearInputKeys().
// #ifndef IMGUI_DISABLE_OBSOLETE_FUNCTIONS
//-----------------------------------------------------------------------------
// [SECTION] Misc data structures (ImGuiInputTextCallbackData, ImGuiSizeCallbackData, ImGuiPayload)
//-----------------------------------------------------------------------------
// Shared state of InputText(), passed as an argument to your callback when a InputTextFlags_Callback* flag is used.
// The callback function should return 0 by default.
// Callbacks (follow a flag name and see comments in InputTextFlags_ declarations for more details)
// - InputTextFlags_CallbackEdit:        Callback on buffer edit. Note that InputText() already returns true on edit + you can always use IsItemEdited(). The callback is useful to manipulate the underlying buffer while focus is active.
// - InputTextFlags_CallbackAlways:      Callback on each iteration
// - InputTextFlags_CallbackCompletion:  Callback on pressing TAB
// - InputTextFlags_CallbackHistory:     Callback on pressing Up/Down arrows
// - InputTextFlags_CallbackCharFilter:  Callback on character inputs to replace or discard them. Modify 'EventChar' to replace or discard, or return 1 in callback to discard.
// - InputTextFlags_CallbackResize:      Callback on buffer capacity changes request (beyond 'buf_size' parameter value), allowing the string to grow.
struct ImGuiInputTextCallbackData { 
	ctx &C.ImGuiContext
// Parent UI context
	eventFlag InputTextFlags
// One InputTextFlags_Callback*    // Read-only
	flags InputTextFlags
// What user passed to InputText()      // Read-only
	userData voidptr
// What user passed to InputText()      // Read-only
// Arguments for the different callback events
// - During Resize callback, Buf will be same as your input buffer.
// - However, during Completion/History/Always callback, Buf always points to our own internal data (it is not the same as your buffer)! Changes to it will be reflected into your own buffer shortly after the callback.
// - To modify the text buffer in a callback, prefer using the InsertChars() / DeleteChars() function. InsertChars() will take care of calling the resize callback if necessary.
// - If you know your edits are not going to resize the underlying buffer allocation, you may modify the contents of 'Buf[]' directly. You need to update 'BufTextLen' accordingly (0 <= BufTextLen < BufSize) and set 'BufDirty'' to true so InputText can update its internal state.
	eventChar C.ImWchar
// Character input                      // Read-write   // [CharFilter] Replace character with another one, or set to zero to drop. return 1 is equivalent to setting EventChar=0;
	eventKey Key
// Key pressed (Up/Down/TAB)            // Read-only    // [Completion,History]
	buf &i8
// Text buffer                          // Read-write   // [Resize] Can replace pointer / [Completion,History,Always] Only write to pointed data, don't replace the actual pointer!
	bufTextLen int
// Text length (in bytes)               // Read-write   // [Resize,Completion,History,Always] Exclude zero-terminator storage. In C land: == strlen(some_text), in C++ land: string.length()
	bufSize int
// Buffer size (in bytes) = capacity+1  // Read-only    // [Resize,Completion,History,Always] Include zero-terminator storage. In C land == ARRAYSIZE(my_char_array), in C++ land: string.capacity()+1
	bufDirty bool
// Set if you modify Buf/BufTextLen!    // Write        // [Completion,History,Always]
	cursorPos int
//                                      // Read-write   // [Completion,History,Always]
	selectionStart int
//                                      // Read-write   // [Completion,History,Always] == to SelectionEnd when no selection)
	selectionEnd int
}
@[c:'ImGuiInputTextCallbackData_DeleteChars']
fn input_text_callback_data_delete_chars(self &ImGuiInputTextCallbackData, pos int, bytes_count int)

@[c:'ImGuiInputTextCallbackData_InsertChars']
fn input_text_callback_data_insert_chars(self &ImGuiInputTextCallbackData, pos int, text &i8, text_end &i8)

@[c:'ImGuiInputTextCallbackData_SelectAll']
fn input_text_callback_data_select_all(self &ImGuiInputTextCallbackData)

@[c:'ImGuiInputTextCallbackData_ClearSelection']
fn input_text_callback_data_clear_selection(self &ImGuiInputTextCallbackData)

@[c:'ImGuiInputTextCallbackData_HasSelection']
fn input_text_callback_data_has_selection(self &ImGuiInputTextCallbackData) bool

// Resizing callback data to apply custom constraint. As enabled by SetNextWindowSizeConstraints(). Callback is called during the next Begin().
// NB: For basic min/max size constraint on each axis you don't need to use the callback! The SetNextWindowSizeConstraints() parameters are enough.
struct ImGuiSizeCallbackData { 
	userData voidptr
// Read-only.   What user passed to SetNextWindowSizeConstraints(). Generally store an integer or float in here (need reinterpret_cast<>).
	pos ImVec2
// Read-only.   Window position, for reference.
	currentSize ImVec2
// Read-only.   Current window size.
	desiredSize ImVec2
}
// Data payload for Drag and Drop operations: AcceptDragDropPayload(), GetDragDropPayload()
struct ImGuiPayload { 
// Members
	data voidptr
// Data (copied and owned by dear imgui)
	dataSize int
// Data size
// [Internal]
	sourceId ID
// Source item id
	sourceParentId ID
// Source parent id (if available)
	dataFrameCount int
// Data timestamp
	dataType [33]i8
// Data type tag (short user-supplied string, 32 characters max)
	preview bool
// Set when AcceptDragDropPayload() was called and mouse has been hovering the target item (nb: handle overlapping drag targets)
	delivery bool
}
@[c:'ImGuiPayload_Clear']
fn payload_clear(self &ImGuiPayload)

@[c:'ImGuiPayload_IsDataType']
fn payload_is_data_type(self &ImGuiPayload, type_ &i8) bool

@[c:'ImGuiPayload_IsPreview']
fn payload_is_preview(self &ImGuiPayload) bool

@[c:'ImGuiPayload_IsDelivery']
fn payload_is_delivery(self &ImGuiPayload) bool

//-----------------------------------------------------------------------------
// [SECTION] Helpers  OnceUponAFrame, ImGuiTextFilter, ImGuiTextBuffer, ImGuiStorage, ImGuiListClipper, Math Operators, ImColor)
//-----------------------------------------------------------------------------
// Helper: Unicode defines
// Invalid Unicode code point (standard value).
// Maximum Unicode code point supported by this build.
// Maximum Unicode code point supported by this build.
// #ifdef IMGUI_USE_WCHAR32
// [Internal]
struct ImGuiTextFilter_ImGuiTextRange { 
	b &i8
	e &i8
}
@[c:'ImGuiTextFilter_ImGuiTextRange_empty']
fn text_filter_im_gui_text_range_empty(self &ImGuiTextFilter_ImGuiTextRange) bool

@[c:'ImGuiTextFilter_ImGuiTextRange_split']
fn text_filter_im_gui_text_range_split(self &ImGuiTextFilter_ImGuiTextRange, separator i8, out &ImVector_ImGuiTextFilter_ImGuiTextRange)

// Helper: Parse and apply text filters. In format "aaaaa[,bbbb][,ccccc]"
struct ImGuiTextFilter { 
	inputBuf [256]i8
	filters ImVector_ImGuiTextFilter_ImGuiTextRange
	countGrep int
}
@[c:'ImGuiTextFilter_Draw']
fn text_filter_draw(self &ImGuiTextFilter, label &i8, width f32) bool

// Helper calling InputText+Build
@[c:'ImGuiTextFilter_PassFilter']
fn text_filter_pass_filter(self &ImGuiTextFilter, text &i8, text_end &i8) bool

@[c:'ImGuiTextFilter_Build']
fn text_filter_build(self &ImGuiTextFilter)

@[c:'ImGuiTextFilter_Clear']
fn text_filter_clear(self &ImGuiTextFilter)

@[c:'ImGuiTextFilter_IsActive']
fn text_filter_is_active(self &ImGuiTextFilter) bool

// Helper: Growable text buffer for logging/accumulating text
// (this could be called 'ImGuiTextBuilder' / 'ImGuiStringBuilder')
struct ImGuiTextBuffer { 
	buf ImVector_char
}
@[c:'ImGuiTextBuffer_begin']
fn text_buffer_begin(self &ImGuiTextBuffer) &i8

@[c:'ImGuiTextBuffer_end']
fn text_buffer_end(self &ImGuiTextBuffer) &i8

// Buf is zero-terminated, so end() will point on the zero-terminator
@[c:'ImGuiTextBuffer_size']
fn text_buffer_size(self &ImGuiTextBuffer) int

@[c:'ImGuiTextBuffer_empty']
fn text_buffer_empty(self &ImGuiTextBuffer) bool

@[c:'ImGuiTextBuffer_clear']
fn text_buffer_clear(self &ImGuiTextBuffer)

@[c:'ImGuiTextBuffer_resize']
fn text_buffer_resize(self &ImGuiTextBuffer, size int)

// Similar to resize(0) on ImVector: empty string but don't free buffer.
@[c:'ImGuiTextBuffer_reserve']
fn text_buffer_reserve(self &ImGuiTextBuffer, capacity int)

@[c:'ImGuiTextBuffer_c_str']
fn text_buffer_c_str(self &ImGuiTextBuffer) &i8

@[c:'ImGuiTextBuffer_append']
fn text_buffer_append(self &ImGuiTextBuffer, str &i8, str_end &i8)

@[c2v_variadic]
@[c:'ImGuiTextBuffer_appendf']
fn text_buffer_appendf(self &ImGuiTextBuffer, fmt &i8)

@[c:'ImGuiTextBuffer_appendfv']
fn text_buffer_appendfv(self &ImGuiTextBuffer, fmt &i8, args C.va_list)

// [Internal] Key+Value for ImGuiStorage
struct ImGuiStoragePair { 
	key ID
}
// Helper: Key->Value storage
// Typically you don't have to worry about this since a storage is held within each Window.
// We use it to e.g. store collapse state for a tree (Int 0/1)
// This is optimized for efficient lookup (dichotomy into a contiguous buffer) and rare insertion (typically tied to user interactions aka max once a frame)
// You can use it as custom user storage for temporary values. Declare your own storage if, for example:
// - You want to manipulate the open/close state of a particular sub-tree in your interface (tree node uses Int 0/1 to store their state).
// - You want to store custom debug data easily without adding or editing structures in your code (probably not efficient, but convenient)
// Types are NOT stored, so it is up to you to make sure your Key don't collide with different types.
struct ImGuiStorage { 
// [Internal]
	data ImVector_ImGuiStoragePair
}
// - Get***() functions find pair, never add/allocate. Pairs are sorted so a query is O(log N)
// - Set***() functions find pair, insertion on demand if missing.
// - Sorted insertion is costly, paid once. A typical frame shouldn't need to insert any new pair.
@[c:'ImGuiStorage_Clear']
fn storage_clear(self &ImGuiStorage)

@[c:'ImGuiStorage_GetInt']
fn storage_get_int(self &ImGuiStorage, key ID, default_val int) int

@[c:'ImGuiStorage_SetInt']
fn storage_set_int(self &ImGuiStorage, key ID, val int)

@[c:'ImGuiStorage_GetBool']
fn storage_get_bool(self &ImGuiStorage, key ID, default_val bool) bool

@[c:'ImGuiStorage_SetBool']
fn storage_set_bool(self &ImGuiStorage, key ID, val bool)

@[c:'ImGuiStorage_GetFloat']
fn storage_get_float(self &ImGuiStorage, key ID, default_val f32) f32

@[c:'ImGuiStorage_SetFloat']
fn storage_set_float(self &ImGuiStorage, key ID, val f32)

@[c:'ImGuiStorage_GetVoidPtr']
fn storage_get_void_ptr(self &ImGuiStorage, key ID) voidptr

// default_val is NULL
@[c:'ImGuiStorage_SetVoidPtr']
fn storage_set_void_ptr(self &ImGuiStorage, key ID, val voidptr)

// - Get***Ref() functions finds pair, insert on demand if missing, return pointer. Useful if you intend to do Get+Set.
// - References are only valid until a new value is added to the storage. Calling a Set***() function or a Get***Ref() function invalidates the pointer.
// - A typical use case where this is convenient for quick hacking (e.g. add storage during a live Edit&Continue session if you can't modify existing struct)
//      float* pvar = ImGui::GetFloatRef(key); ImGui::SliderFloat("var", pvar, 0, 100.0f); some_var += *pvar;
@[c:'ImGuiStorage_GetIntRef']
fn storage_get_int_ref(self &ImGuiStorage, key ID, default_val int) &int

@[c:'ImGuiStorage_GetBoolRef']
fn storage_get_bool_ref(self &ImGuiStorage, key ID, default_val bool) &bool

@[c:'ImGuiStorage_GetFloatRef']
fn storage_get_float_ref(self &ImGuiStorage, key ID, default_val f32) &f32

@[c:'ImGuiStorage_GetVoidPtrRef']
fn storage_get_void_ptr_ref(self &ImGuiStorage, key ID, default_val voidptr) &voidptr

// Advanced: for quicker full rebuild of a storage (instead of an incremental one), you may add all your contents and then sort once.
@[c:'ImGuiStorage_BuildSortByKey']
fn storage_build_sort_by_key(self &ImGuiStorage)

// Obsolete: use on your own storage if you know only integer are being stored (open/close all tree nodes)
@[c:'ImGuiStorage_SetAllInt']
fn storage_set_all_int(self &ImGuiStorage, val int)

// Helper: Manually clip large list of items.
// If you have lots evenly spaced items and you have random access to the list, you can perform coarse
// clipping based on visibility to only submit items that are in view.
// The clipper calculates the range of visible items and advance the cursor to compensate for the non-visible items we have skipped.
// (Dear ImGui already clip items based on their bounds but: it needs to first layout the item to do so, and generally
//  fetching/submitting your own data incurs additional cost. Coarse clipping using ImGuiListClipper allows you to easily
//  scale using lists with tens of thousands of items without a problem)
// Usage:
//   ImGuiListClipper clipper;
//   clipper.Begin(1000);         // We have 1000 elements, evenly spaced.
//   while (clipper.Step())
//       for (int i = clipper.DisplayStart; i < clipper.DisplayEnd; i++)
//           ImGui::Text("line number %d", i);
// Generally what happens is:
// - Clipper lets you process the first element (DisplayStart = 0, DisplayEnd = 1) regardless of it being visible or not.
// - User code submit that one element.
// - Clipper can measure the height of the first element
// - Clipper calculate the actual range of elements to display based on the current clipping rectangle, position the cursor before the first visible element.
// - User code submit visible elements.
// - The clipper also handles various subtleties related to keyboard/gamepad navigation, wrapping etc.
struct ImGuiListClipper { 
	ctx &C.ImGuiContext
// Parent UI context
	displayStart int
// First item to display, updated by each call to Step()
	displayEnd int
// End of items to display (exclusive)
	itemsCount int
// [Internal] Number of items
	itemsHeight f32
// [Internal] Height of item after a first step and item submission can calculate it
	startPosY f32
// [Internal] Cursor position at the time of Begin() or after table frozen rows are all processed
	startSeekOffsetY f64
// [Internal] Account for frozen rows in a table and initial loss of precision in very large windows.
	tempData voidptr
}
@[c:'ImGuiListClipper_Begin']
fn list_clipper_begin(self &ImGuiListClipper, items_count int, items_height f32)

@[c:'ImGuiListClipper_End']
fn list_clipper_end(self &ImGuiListClipper)

// Automatically called on the last call of Step() that returns false.
@[c:'ImGuiListClipper_Step']
fn list_clipper_step(self &ImGuiListClipper) bool

// Call until it returns false. The DisplayStart/DisplayEnd fields will be set and you can process/draw those items.
// Call IncludeItemByIndex() or IncludeItemsByIndex() *BEFORE* first call to Step() if you need a range of items to not be clipped, regardless of their visibility.
// (Due to alignment / padding of certain items it is possible that an extra item may be included on either end of the display range).
@[c:'ImGuiListClipper_IncludeItemByIndex']
fn list_clipper_include_item_by_index(self &ImGuiListClipper, item_index int)

@[c:'ImGuiListClipper_IncludeItemsByIndex']
fn list_clipper_include_items_by_index(self &ImGuiListClipper, item_begin int, item_end int)

// item_end is exclusive e.g. use (42, 42+1) to make item 42 never clipped.
// Seek cursor toward given item. This is automatically called while stepping.
// - The only reason to call this is: you can use ImGuiListClipper::Begin(INT_MAX) if you don't know item count ahead of time.
// - In this case, after all steps are done, you'll want to call SeekCursorForItem(item_count).
@[c:'ImGuiListClipper_SeekCursorForItem']
fn list_clipper_seek_cursor_for_item(self &ImGuiListClipper, item_index int)

@[c:'ImGuiListClipper_IncludeRangeByIndices']
fn list_clipper_include_range_by_indices(self &ImGuiListClipper, item_begin int, item_end int)

// [renamed in 1.89.9]
@[c:'ImGuiListClipper_ForceDisplayRangeByIndices']
fn list_clipper_force_display_range_by_indices(self &ImGuiListClipper, item_begin int, item_end int)

// [renamed in 1.89.6]
// #ifndef IMGUI_DISABLE_OBSOLETE_FUNCTIONS
// Helpers: ImVec2/C.ImVec4 operators
// - It is important that we are keeping those disabled by default so they don't leak in user space.
// - This is in order to allow user enabling implicit cast operators between ImVec2/C.ImVec4 and their own types (using IM_VEC2_CLASS_EXTRA in imconfig.h)
// - Add '#define IMGUI_DEFINE_MATH_OPERATORS' before including this file (or in imconfig.h) to access courtesy maths operators for ImVec2 and C.ImVec4.
// - We intentionally provide ImVec2*float but not float*ImVec2: this is rare enough and we want to reduce the surface for possible user mistake.
// #ifdef IMGUI_DEFINE_MATH_OPERATORS
// Helpers macros to generate 32-bit encoded colors
// - User can declare their own format by #defining the 5 _SHIFT/_MASK macros in their imconfig file.
// - Any setting other than the default will need custom backend support. The only standard backend that supports anything else than the default is DirectX9.
// #ifdef IMGUI_USE_BGRA_PACKED_COLOR
// #ifndef IM_COL32_R_SHIFT
// Opaque white = 0xFFFFFFFF
// Opaque black
// Transparent black = 0x00000000
// Helper: ImColor() implicitly converts colors to either ImU32 (packed 4x1 byte) or C.ImVec4 (4x1 float)
// Prefer using IM_COL32() macros if you want a guaranteed compile-time ImU32 for usage with ImDrawList API.
// **Avoid storing ImColor! Store either u32 of C.ImVec4. This is not a full-featured color class. MAY OBSOLETE.
// **None of the ImGui API are using ImColor directly but you can use it as a convenience to pass colors in either ImU32 or C.ImVec4 formats. Explicitly cast to ImU32 or C.ImVec4 if needed.
struct ImColor { 
	value C.ImVec4
}
// FIXME-OBSOLETE: May need to obsolete/cleanup those helpers.
@[c:'ImColor_SetHSV']
fn im_color_set_hsv(self &ImColor, h f32, s f32, v f32, a f32)

@[c:'ImColor_HSV']
fn im_color_hsv(h f32, s f32, v f32, a f32) ImColor

//-----------------------------------------------------------------------------
// [SECTION] Multi-Select API flags and structures  MultiSelectFlags, ImGuiSelectionRequestType, ImGuiSelectionRequest, ImGuiMultiSelectIO, ImGuiSelectionBasicStorage)
//-----------------------------------------------------------------------------
// Multi-selection system
// Documentation at: https://github.com/ocornut/imgui/wiki/Multi-Select
// - Refer to 'Demo->Widgets->Selection State & Multi-Select' for demos using this.
// - This system implements standard multi-selection idioms (CTRL+Mouse/Keyboard, SHIFT+Mouse/Keyboard, etc)
//   with support for clipper (skipping non-visible items), box-select and many other details.
// - Selectable(), Checkbox() are supported but custom widgets may use it as well.
// - TreeNode() is technically supported but... using this correctly is more complicated: you need some sort of linear/random access to your tree,
//   which is suited to advanced trees setups also implementing filters and clipper. We will work toward simplifying and demoing it.
// - In the spirit of Dear ImGui design, your code owns actual selection data.
//   This is designed to allow all kinds of selection storage you may use in your application e.g. set/map/hash.
// About ImGuiSelectionBasicStorage:
// - This is an optional helper to store a selection state and apply selection requests.
// - It is used by our demos and provided as a convenience to quickly implement multi-selection.
// Usage:
// - Identify submitted items with SetNextItemSelectionUserData(), most likely using an index into your current data-set.
// - Store and maintain actual selection data using persistent object identifiers.
// - Usage flow:
//     BEGIN - (1) Call BeginMultiSelect() and retrieve the ImGuiMultiSelectIO* result.
//           - (2) Honor request list (SetAll/SetRange requests) by updating your selection data. Same code as Step 6.
//           - (3) [If using clipper] You need to make sure RangeSrcItem is always submitted. Calculate its index and pass to clipper.IncludeItemByIndex(). If storing indices in SelectionUserData, a simple clipper.IncludeItemByIndex(ms_io->RangeSrcItem) call will work.
//     LOOP  - (4) Submit your items with SetNextItemSelectionUserData() + Selectable()/TreeNode() calls.
//     END   - (5) Call EndMultiSelect() and retrieve the ImGuiMultiSelectIO* result.
//           - (6) Honor request list (SetAll/SetRange requests) by updating your selection data. Same code as Step 2.
//     If you submit all items (no clipper), Step 2 and 3 are optional and will be handled by each item themselves. It is fine to always honor those steps.
// About SelectionUserData:
// - This can store an application-defined identifier (e.g. index or pointer) submitted via SetNextItemSelectionUserData().
// - In return we store them into RangeSrcItem/RangeFirstItem/RangeLastItem and other fields in ImGuiMultiSelectIO.
// - Most applications will store an object INDEX, hence the chosen name and type. Storing an index is natural, because
//   SetRange requests will give you two end-points and you will need to iterate/interpolate between them to update your selection.
// - However it is perfectly possible to store a POINTER or another IDENTIFIER inside SelectionUserData.
//   Our system never assume that you identify items by indices, it never attempts to interpolate between two values.
// - If you enable MultiSelectFlags_NoRangeSelect then it is guaranteed that you will never have to interpolate
//   between two SelectionUserData, which may be a convenient way to use part of the feature with less code work.
// - As most users will want to store an index, for convenience and to reduce confusion we use ImS64 instead of void*,
//   being syntactically easier to downcast. Feel free to reinterpret_cast and store a pointer inside.
// Flags for BeginMultiSelect()
enum MultiSelectFlags_ {
 none = 0
 single_select = 1 << 0
// Disable selecting more than one item. This is available to allow single-selection code to share same code/logic if desired. It essentially disables the main purpose of BeginMultiSelect() tho!
 no_select_all = 1 << 1
// Disable CTRL+A shortcut to select all.
 no_range_select = 1 << 2
// Disable Shift+selection mouse/keyboard support (useful for unordered 2D selection). With BoxSelect is also ensure contiguous SetRange requests are not combined into one. This allows not handling interpolation in SetRange requests.
 no_auto_select = 1 << 3
// Disable selecting items when navigating (useful for e.g. supporting range-select in a list of checkboxes).
 no_auto_clear = 1 << 4
// Disable clearing selection when navigating or selecting another one (generally used with MultiSelectFlags_NoAutoSelect. useful for e.g. supporting range-select in a list of checkboxes).
 no_auto_clear_on_reselect = 1 << 5
// Disable clearing selection when clicking/selecting an already selected item.
 box_select1d = 1 << 6
// Enable box-selection with same width and same x pos items (e.g. full row Selectable()). Box-selection works better with little bit of spacing between items hit-box in order to be able to aim at empty space.
 box_select2d = 1 << 7
// Enable box-selection with varying width or varying x pos items support (e.g. different width labels, or 2D layout/grid). This is slower: alters clipping logic so that e.g. horizontal movements will update selection of normally clipped items.
 box_select_no_scroll = 1 << 8
// Disable scrolling when box-selecting near edges of scope.
 clear_on_escape = 1 << 9
// Clear selection when pressing Escape while scope is focused.
 clear_on_click_void = 1 << 10
// Clear selection when clicking on empty location within scope.
 scope_window = 1 << 11
// Scope for _BoxSelect and _ClearOnClickVoid is whole window (Default). Use if BeginMultiSelect() covers a whole window or used a single time in same window.
 scope_rect = 1 << 12
// Scope for _BoxSelect and _ClearOnClickVoid is rectangle encompassing BeginMultiSelect()/EndMultiSelect(). Use if BeginMultiSelect() is called multiple times in same window.
 select_on_click = 1 << 13
// Apply selection on mouse down when clicking on unselected item. (Default)
 select_on_click_release = 1 << 14
// Apply selection on mouse release when clicking an unselected item. Allow dragging an unselected item without altering selection.
//ImGuiMultiSelectFlags_RangeSelect2d       = 1 << 15,  // Shift+Selection uses 2d geometry instead of linear sequence, so possible to use Shift+up/down to select vertically in grid. Analogous to what BoxSelect does.
 nav_wrap_x = 1 << 16
}

// Main IO structure returned by BeginMultiSelect()/EndMultiSelect().
// This mainly contains a list of selection requests.
// - Use 'Demo->Tools->Debug Log->Selection' to see requests as they happen.
// - Some fields are only useful if your list is dynamic and allows deletion (getting post-deletion focus/state right is shown in the demo)
// - Below: who reads/writes each fields? 'r'=read, 'w'=write, 'ms'=multi-select code, 'app'=application/user code.
struct ImGuiMultiSelectIO { 
//------------------------------------------// BeginMultiSelect / EndMultiSelect
	requests ImVector_ImGuiSelectionRequest
//  ms:w, app:r     /  ms:w  app:r   // Requests to apply to your selection data.
	rangeSrcItem SelectionUserData
//  ms:w  app:r     /                // (If using clipper) Begin: Source item (often the first selected item) must never be clipped: use clipper.IncludeItemByIndex() to ensure it is submitted.
	navIdItem SelectionUserData
//  ms:w, app:r     /                // (If using deletion) Last known SetNextItemSelectionUserData() value for NavId (if part of submitted items).
	navIdSelected bool
//  ms:w, app:r     /        app:r   // (If using deletion) Last known selection state for NavId (if part of submitted items).
	rangeSrcReset bool
//        app:w     /  ms:r          // (If using deletion) Set before EndMultiSelect() to reset ResetSrcItem (e.g. if deleted selection).
	itemsCount int
}
// Selection request type
enum ImGuiSelectionRequestType {
 selection_request_type_none = 0
 selection_request_type_set_all
// Request app to clear selection (if Selected==false) or select all items (if Selected==true). We cannot set RangeFirstItem/RangeLastItem as its contents is entirely up to user (not necessarily an index)
 selection_request_type_set_range
}

// Selection request item
struct ImGuiSelectionRequest { 
//------------------------------------------// BeginMultiSelect / EndMultiSelect
	type ImGuiSelectionRequestType
//  ms:w, app:r     /  ms:w, app:r   // Request type. You'll most often receive 1 Clear + 1 SetRange with a single-item range.
	selected bool
//  ms:w, app:r     /  ms:w, app:r   // Parameter for SetAll/SetRange requests (true = select, false = unselect)
	rangeDirection ImS8
//                  /  ms:w  app:r   // Parameter for SetRange request: +1 when RangeFirstItem comes before RangeLastItem, -1 otherwise. Useful if you want to preserve selection order on a backward Shift+Click.
	rangeFirstItem SelectionUserData
//                  /  ms:w, app:r   // Parameter for SetRange request (this is generally == RangeSrcItem when shift selecting from top to bottom).
	rangeLastItem SelectionUserData
}
// Optional helper to store multi-selection state + apply multi-selection requests.
// - Used by our demos and provided as a convenience to easily implement basic multi-selection.
// - Iterate selection with 'void* it = NULL; ID id; while (selection.GetNextSelectedItem(&it, &id)) { ... }'
//   Or you can check 'if (Contains(id)) { ... }' for each possible object if their number is not too high to iterate.
// - USING THIS IS NOT MANDATORY. This is only a helper and not a required API.
// To store a multi-selection, in your application you could:
// - Use this helper as a convenience. We use our simple key->value ImGuiStorage as a std::set ID> replacement.
// - Use your own external storage: e.g. std::set<MyObjectId>, std::vector<MyObjectId>, interval trees, intrusively stored selection etc.
// In ImGuiSelectionBasicStorage we:
// - always use indices in the multi-selection API (passed to SetNextItemSelectionUserData(), retrieved in ImGuiMultiSelectIO)
// - use the AdapterIndexToStorageId() indirection layer to abstract how persistent selection data is derived from an index.
// - use decently optimized logic to allow queries and insertion of very large selection sets.
// - do not preserve selection order.
// Many combinations are possible depending on how you prefer to store your items and how you prefer to store your selection.
// Large applications are likely to eventually want to get rid of this indirection layer and do their own thing.
// See https://github.com/ocornut/imgui/wiki/Multi-Select for details and pseudo-code using this helper.
struct ImGuiSelectionBasicStorage { 
// Members
	size int
//          // Number of selected items, maintained by this helper.
	preserveOrder bool
// = false  // GetNextSelectedItem() will return ordered selection (currently implemented by two additional sorts of selection. Could be improved)
	userData voidptr
// = NULL   // User data for use by adapter function        // e.g. selection.UserData = (void*)my_items;
	adapterIndexToStorageId fn (&ImGuiSelectionBasicStorage, int) ID
// e.g. selection.AdapterIndexToStorageId = [](ImGuiSelectionBasicStorage* self, int idx) { return ((MyItems**)self->UserData)[idx]->ID; };
	_SelectionOrder int
// [Internal] Increasing counter to store selection order
	_Storage ImGuiStorage
}
@[c:'ImGuiSelectionBasicStorage_ApplyRequests']
fn selection_basic_storage_apply_requests(self &ImGuiSelectionBasicStorage, ms_io &ImGuiMultiSelectIO)

// Apply selection requests coming from BeginMultiSelect() and EndMultiSelect() functions. It uses 'items_count' passed to BeginMultiSelect()
@[c:'ImGuiSelectionBasicStorage_Contains']
fn selection_basic_storage_contains(self &ImGuiSelectionBasicStorage, id ID) bool

// Query if an item id is in selection.
@[c:'ImGuiSelectionBasicStorage_Clear']
fn selection_basic_storage_clear(self &ImGuiSelectionBasicStorage)

// Clear selection
@[c:'ImGuiSelectionBasicStorage_Swap']
fn selection_basic_storage_swap(self &ImGuiSelectionBasicStorage, r &ImGuiSelectionBasicStorage)

// Swap two selections
@[c:'ImGuiSelectionBasicStorage_SetItemSelected']
fn selection_basic_storage_set_item_selected(self &ImGuiSelectionBasicStorage, id ID, selected bool)

// Add/remove an item from selection (generally done by ApplyRequests() function)
@[c:'ImGuiSelectionBasicStorage_GetNextSelectedItem']
fn selection_basic_storage_get_next_selected_item(self &ImGuiSelectionBasicStorage, opaque_it &voidptr, out_id  ID) bool

// Iterate selection with 'void* it = NULL; ID id; while (selection.GetNextSelectedItem(&it, &id)) { ... }'
@[c:'ImGuiSelectionBasicStorage_GetStorageIdFromIndex']
fn selection_basic_storage_get_storage_id_from_index(self &ImGuiSelectionBasicStorage, idx int) ID

// Convert index to item id based on provided adapter.
// Optional helper to apply multi-selection requests to existing randomly accessible storage.
// Convenient if you want to quickly wire multi-select API on e.g. an array of bool or items storing their own selection state.
struct ImGuiSelectionExternalStorage { 
// Members
	userData voidptr
// User data for use by adapter function                                // e.g. selection.UserData = (void*)my_items;
	adapterSetItemSelected fn (&ImGuiSelectionExternalStorage, int, bool)
}
@[c:'ImGuiSelectionExternalStorage_ApplyRequests']
fn selection_external_storage_apply_requests(self &ImGuiSelectionExternalStorage, ms_io &ImGuiMultiSelectIO)

// Apply selection requests by using AdapterSetItemSelected() calls
//-----------------------------------------------------------------------------
// [SECTION] Drawing API (ImDrawCmd, ImDrawIdx, ImDrawVert, ImDrawChannel, ImDrawListSplitter, ImDrawListFlags, ImDrawList, ImDrawData)
// Hold a series of drawing commands. The user provides a renderer for ImDrawData which essentially contains an array of ImDrawList.
//-----------------------------------------------------------------------------
// The maximum line width to bake anti-aliased textures for. Build atlas with ImFontAtlasFlags_NoBakedLines to disable baking.
// #ifndef IM_DRAWLIST_TEX_LINES_WIDTH_MAX
// ImDrawCallback: Draw callbacks for advanced uses [configurable type: override in imconfig.h]
// NB: You most likely do NOT need to use draw callbacks just to create your own widget or customized UI rendering,
// you can poke into the draw list for that! Draw callback may be useful for example to:
//  A) Change your GPU render state,
//  B) render a complex 3D scene inside a UI element without an intermediate texture/render target, etc.
// The expected behavior from your rendering function is 'if (cmd.UserCallback != NULL) { cmd.UserCallback(parent_list, cmd); } else { RenderTriangles() }'
// If you want to override the signature of ImDrawCallback, you can simply use e.g. '#define ImDrawCallback MyDrawCallback' (in imconfig.h) + update rendering backend accordingly.
type ImDrawCallback = fn (&ImDrawList, &ImDrawCmd)
// #ifndef ImDrawCallback
// Special Draw callback value to request renderer backend to reset the graphics/render state.
// The renderer backend needs to handle this special value, otherwise it will crash trying to call a function at this address.
// This is useful, for example, if you submitted callbacks which you know have altered the render state and you want it to be restored.
// Render state is not reset by default because they are many perfectly useful way of altering render state (e.g. changing shader/blending settings before an Image call).
// Typically, 1 command = 1 GPU draw call (unless command is a callback)
// - VtxOffset: When 'io.BackendFlags & BackendFlags_RendererHasVtxOffset' is enabled,
//   this fields allow us to render meshes larger than 64K vertices while keeping 16-bit indices.
//   Backends made for <1.71. will typically ignore the VtxOffset fields.
// - The ClipRect/TextureId/VtxOffset fields must be contiguous as we memcmp() them together (this is asserted for).
struct ImDrawCmd { 
	clipRect C.ImVec4
// 4*4  // Clipping rectangle (x1, y1, x2, y2). Subtract ImDrawData->DisplayPos to get clipping rectangle in "viewport" coordinates
	textureId ImTextureID
// 4-8  // User-provided texture ID. Set by user in ImfontAtlas::SetTexID() for fonts or passed to Image*() functions. Ignore if never using images or multiple fonts atlas.
	vtxOffset u32
// 4    // Start offset in vertex buffer. BackendFlags_RendererHasVtxOffset: always 0, otherwise may be >0 to support meshes larger than 64K vertices with 16-bit indices.
	idxOffset u32
// 4    // Start offset in index buffer.
	elemCount u32
// 4    // Number of indices (multiple of 3) to be rendered as triangles. Vertices are stored in the callee ImDrawList's vtx_buffer[] array, indices in idx_buffer[].
	userCallback ImDrawCallback
// 4-8  // If != NULL, call the function instead of rendering the vertices. clip_rect and texture_id will be set normally.
	userCallbackData voidptr
// 4-8  // Callback user data (when UserCallback != NULL). If called AddCallback() with size == 0, this is a copy of the AddCallback() argument. If called AddCallback() with size > 0, this is pointing to a buffer where data is stored.
	userCallbackDataSize int
// 4 // Size of callback user data when using storage, otherwise 0.
	userCallbackDataOffset int
}
// Since 1.83: returns ImTextureID associated with this draw call. Warning: DO NOT assume this is always same as 'TextureId' (we will change this function for an upcoming feature)
@[c:'ImDrawCmd_GetTexID']
fn im_draw_cmd_get_tex_id(self &ImDrawCmd) ImTextureID

// Vertex layout
struct ImDrawVert { 
	pos ImVec2
	uv ImVec2
	col ImU32
}
// You can override the vertex format layout by defining IMGUI_OVERRIDE_DRAWVERT_STRUCT_LAYOUT in imconfig.h
// The code expect ImVec2 pos (8 bytes), ImVec2 uv (8 bytes), ImU32 col (4 bytes), but you can re-order them or add other fields as needed to simplify integration in your engine.
// The type has to be described within the macro (you can either declare the struct or use a typedef). This is because ImVec2/ImU32 are likely not declared at the time you'd want to set your type up.
// NOTE: IMGUI DOESN'T CLEAR THE STRUCTURE AND DOESN'T CALL A CONSTRUCTOR SO ANY CUSTOM FIELD WILL BE UNINITIALIZED. IF YOU ADD EXTRA FIELDS (SUCH AS A 'Z' COORDINATES) YOU WILL NEED TO CLEAR THEM DURING RENDER OR TO IGNORE THEM.
// #ifndef IMGUI_OVERRIDE_DRAWVERT_STRUCT_LAYOUT
// [Internal] For use by ImDrawList
struct ImDrawCmdHeader { 
	clipRect C.ImVec4
	textureId ImTextureID
	vtxOffset u32
}
// [Internal] For use by ImDrawListSplitter
struct ImDrawChannel { 
	_CmdBuffer ImVector_ImDrawCmd
	_IdxBuffer ImVector_ImDrawIdx
}
// Split/Merge functions are used to split the draw list into different layers which can be drawn into out of order.
// This is used by the Columns/Tables API, so items of each column can be batched together in a same draw call.
struct ImDrawListSplitter { 
	_Current int
// Current channel number (0)
	_Count int
// Number of active channels (1+)
	_Channels ImVector_ImDrawChannel
}
@[c:'ImDrawListSplitter_Clear']
fn im_draw_list_splitter_clear(self &ImDrawListSplitter)

// Do not clear Channels[] so our allocations are reused next frame
@[c:'ImDrawListSplitter_ClearFreeMemory']
fn im_draw_list_splitter_clear_free_memory(self &ImDrawListSplitter)

@[c:'ImDrawListSplitter_Split']
fn im_draw_list_splitter_split(self &ImDrawListSplitter, draw_list &ImDrawList, count int)

@[c:'ImDrawListSplitter_Merge']
fn im_draw_list_splitter_merge(self &ImDrawListSplitter, draw_list &ImDrawList)

@[c:'ImDrawListSplitter_SetCurrentChannel']
fn im_draw_list_splitter_set_current_channel(self &ImDrawListSplitter, draw_list &ImDrawList, channel_idx int)

// Flags for ImDrawList functions
// (Legacy: bit 0 must always correspond to ImDrawFlags_Closed to be backward compatible with old API using a bool. Bits 1..3 must be unused)
enum ImDrawFlags_ {
	none = 0
	closed = 1 << 0
// PathStroke(), AddPolyline(): specify that shape should be closed (Important: this is always == 1 for legacy reason)
	round_corners_top_left = 1 << 4
// AddRect(), AddRectFilled(), PathRect(): enable rounding top-left corner only (when rounding > 0.0f, we default to all corners). Was 0x01.
	round_corners_top_right = 1 << 5
// AddRect(), AddRectFilled(), PathRect(): enable rounding top-right corner only (when rounding > 0.0f, we default to all corners). Was 0x02.
	round_corners_bottom_left = 1 << 6
// AddRect(), AddRectFilled(), PathRect(): enable rounding bottom-left corner only (when rounding > 0.0f, we default to all corners). Was 0x04.
	round_corners_bottom_right = 1 << 7
// AddRect(), AddRectFilled(), PathRect(): enable rounding bottom-right corner only (when rounding > 0.0f, we default to all corners). Wax 0x08.
	round_corners_none = 1 << 8
// AddRect(), AddRectFilled(), PathRect(): disable rounding on all corners (when rounding > 0.0f). This is NOT zero, NOT an implicit flag!
	round_corners_top = 1 << 4 | 1 << 5
	round_corners_bottom = 1 << 6 | 1 << 7
	round_corners_left = 1 << 6 | 1 << 4
	round_corners_right = 1 << 7 | 1 << 5
	round_corners_all = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	round_corners_default_ = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
// Default to ALL corners if none of the _RoundCornersXX flags are specified.
	round_corners_mask_ = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8
}

// Flags for ImDrawList instance. Those are set automatically by ImGui:: functions from ImGuiIO settings, and generally not manipulated directly.
// It is however possible to temporarily alter flags between calls to ImDrawList:: functions.
enum ImDrawListFlags_ {
	none = 0
	anti_aliased_lines = 1 << 0
// Enable anti-aliased lines/borders (*2 the number of triangles for 1.0f wide line or lines thin enough to be drawn using textures, otherwise *3 the number of triangles)
	anti_aliased_lines_use_tex = 1 << 1
// Enable anti-aliased lines/borders using textures when possible. Require backend to render with bilinear filtering (NOT point/nearest filtering).
	anti_aliased_fill = 1 << 2
// Enable anti-aliased edge around filled shapes (rounded rectangles, circles).
	allow_vtx_offset = 1 << 3
}

// Draw command list
// This is the low-level list of polygons that ImGui:: functions are filling. At the end of the frame,
// all command lists are passed to your ImGuiIO::RenderDrawListFn function for rendering.
// Each dear imgui window contains its own ImDrawList. You can use ImGui::GetWindowDrawList() to
// access the current window draw list and draw custom primitives.
// You can interleave normal ImGui:: calls and adding primitives to the current draw list.
// In single viewport mode, top-left is == GetMainViewport()->Pos (generally 0,0), bottom-right is == GetMainViewport()->Pos+Size (generally io.DisplaySize).
// You are totally free to apply whatever transformation matrix you want to the data (depending on the use of the transformation you may want to apply it to ClipRect as well!)
// Important: Primitives are always added to the list and not culled (culling is done at higher-level by ImGui:: functions), if you use this API a lot consider coarse culling your drawn objects.
struct ImDrawList { 
// This is what you have to render
	cmdBuffer ImVector_ImDrawCmd
// Draw commands. Typically 1 command = 1 GPU draw call, unless the command is a callback.
	idxBuffer ImVector_ImDrawIdx
// Index buffer. Each command consume ImDrawCmd::ElemCount of those
	vtxBuffer ImVector_ImDrawVert
// Vertex buffer.
	flags ImDrawListFlags
// Flags, you may poke into these to adjust anti-aliasing settings per-primitive.
// [Internal, used while building lists]
	_VtxCurrentIdx u32
// [Internal] generally == VtxBuffer.Size unless we are past 64K vertices, in which case this gets reset to 0.
	_Data &C.ImDrawListSharedData
// Pointer to shared draw data (you can use ImGui::GetDrawListSharedData() to get the one from current ImGui context)
	_VtxWritePtr &ImDrawVert
// [Internal] point within VtxBuffer.Data after each add command (to avoid using the ImVector<> operators too much)
	_IdxWritePtr &ImDrawIdx
// [Internal] point within IdxBuffer.Data after each add command (to avoid using the ImVector<> operators too much)
	_Path ImVector_ImVec2
// [Internal] current path building
	_CmdHeader ImDrawCmdHeader
// [Internal] template of active commands. Fields should match those of CmdBuffer.back().
	_Splitter ImDrawListSplitter
// [Internal] for channels api (note: prefer using your own persistent instance of ImDrawListSplitter!)
	_ClipRectStack ImVector_ImVec4
// [Internal]
	_TextureIdStack ImVector_ImTextureID
// [Internal]
	_CallbacksDataBuf ImVector_ImU8
// [Internal]
	_FringeScale f32
// [Internal] anti-alias fringe is scaled by this value, this helps to keep things sharp while zooming at vertex buffer content
	_OwnerName &i8
// Pointer to owner window's name for debugging
// Obsolete names
//inline  void  AddEllipse(const ImVec2& center, float radius_x, float radius_y, ImU32 col, float rot = 0.0f, int num_segments = 0, float thickness = 1.0f) { AddEllipse(center, ImVec2(radius_x, radius_y), col, rot, num_segments, thickness); } // OBSOLETED in 1.90.5 (Mar 2024)
//inline  void  AddEllipseFilled(const ImVec2& center, float radius_x, float radius_y, ImU32 col, float rot = 0.0f, int num_segments = 0) { AddEllipseFilled(center, ImVec2(radius_x, radius_y), col, rot, num_segments); }                        // OBSOLETED in 1.90.5 (Mar 2024)
//inline  void  PathEllipticalArcTo(const ImVec2& center, float radius_x, float radius_y, float rot, float a_min, float a_max, int num_segments = 0) { PathEllipticalArcTo(center, ImVec2(radius_x, radius_y), rot, a_min, a_max, num_segments); } // OBSOLETED in 1.90.5 (Mar 2024)
//inline  void  AddBezierCurve(const ImVec2& p1, const ImVec2& p2, const ImVec2& p3, const ImVec2& p4, ImU32 col, float thickness, int num_segments = 0) { AddBezierCubic(p1, p2, p3, p4, col, thickness, num_segments); }                         // OBSOLETED in 1.80 (Jan 2021)
}
@[c:'ImDrawList_PushClipRect']
fn im_draw_list_push_clip_rect(self &ImDrawList, clip_rect_min ImVec2, clip_rect_max ImVec2, intersect_with_current_clip_rect bool)

// Render-level scissoring. This is passed down to your render function but not used for CPU-side coarse clipping. Prefer using higher-level ImGui::PushClipRect() to affect logic (hit-testing and widget culling)
@[c:'ImDrawList_PushClipRectFullScreen']
fn im_draw_list_push_clip_rect_full_screen(self &ImDrawList)

@[c:'ImDrawList_PopClipRect']
fn im_draw_list_pop_clip_rect(self &ImDrawList)

@[c:'ImDrawList_PushTextureID']
fn im_draw_list_push_texture_id(self &ImDrawList, texture_id ImTextureID)

@[c:'ImDrawList_PopTextureID']
fn im_draw_list_pop_texture_id(self &ImDrawList)

@[c:'ImDrawList_GetClipRectMin']
fn im_draw_list_get_clip_rect_min(self &ImDrawList) ImVec2

@[c:'ImDrawList_GetClipRectMax']
fn im_draw_list_get_clip_rect_max(self &ImDrawList) ImVec2

// Primitives
// - Filled shapes must always use clockwise winding order. The anti-aliasing fringe depends on it. Counter-clockwise shapes will have "inward" anti-aliasing.
// - For rectangular primitives, "p_min" and "p_max" represent the upper-left and lower-right corners.
// - For circle primitives, use "num_segments == 0" to automatically calculate tessellation (preferred).
//   In older versions (until Dear ImGui 1.77) the AddCircle functions defaulted to num_segments == 12.
//   In future versions we will use textures to provide cheaper and higher-quality circles.
//   Use AddNgon() and AddNgonFilled() functions if you need to guarantee a specific number of sides.
@[c:'ImDrawList_AddLine']
fn im_draw_list_add_line(self &ImDrawList, p1 ImVec2, p2 ImVec2, col ImU32)

// Implied thickness = 1.0f
@[c:'ImDrawList_AddLineEx']
fn im_draw_list_add_line_ex(self &ImDrawList, p1 ImVec2, p2 ImVec2, col ImU32, thickness f32)

@[c:'ImDrawList_AddRect']
fn im_draw_list_add_rect(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32)

// Implied rounding = 0.0f, flags = 0, thickness = 1.0f
@[c:'ImDrawList_AddRectEx']
fn im_draw_list_add_rect_ex(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags, thickness f32)

// a: upper-left, b: lower-right (== upper-left + size)
@[c:'ImDrawList_AddRectFilled']
fn im_draw_list_add_rect_filled(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32)

// Implied rounding = 0.0f, flags = 0
@[c:'ImDrawList_AddRectFilledEx']
fn im_draw_list_add_rect_filled_ex(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags)

// a: upper-left, b: lower-right (== upper-left + size)
@[c:'ImDrawList_AddRectFilledMultiColor']
fn im_draw_list_add_rect_filled_multi_color(self &ImDrawList, p_min ImVec2, p_max ImVec2, col_upr_left ImU32, col_upr_right ImU32, col_bot_right ImU32, col_bot_left ImU32)

@[c:'ImDrawList_AddQuad']
fn im_draw_list_add_quad(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32)

// Implied thickness = 1.0f
@[c:'ImDrawList_AddQuadEx']
fn im_draw_list_add_quad_ex(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32, thickness f32)

@[c:'ImDrawList_AddQuadFilled']
fn im_draw_list_add_quad_filled(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32)

@[c:'ImDrawList_AddTriangle']
fn im_draw_list_add_triangle(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32)

// Implied thickness = 1.0f
@[c:'ImDrawList_AddTriangleEx']
fn im_draw_list_add_triangle_ex(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32, thickness f32)

@[c:'ImDrawList_AddTriangleFilled']
fn im_draw_list_add_triangle_filled(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32)

@[c:'ImDrawList_AddCircle']
fn im_draw_list_add_circle(self &ImDrawList, center ImVec2, radius f32, col ImU32)

// Implied num_segments = 0, thickness = 1.0f
@[c:'ImDrawList_AddCircleEx']
fn im_draw_list_add_circle_ex(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int, thickness f32)

@[c:'ImDrawList_AddCircleFilled']
fn im_draw_list_add_circle_filled(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

@[c:'ImDrawList_AddNgon']
fn im_draw_list_add_ngon(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

// Implied thickness = 1.0f
@[c:'ImDrawList_AddNgonEx']
fn im_draw_list_add_ngon_ex(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int, thickness f32)

@[c:'ImDrawList_AddNgonFilled']
fn im_draw_list_add_ngon_filled(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

@[c:'ImDrawList_AddEllipse']
fn im_draw_list_add_ellipse(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32)

// Implied rot = 0.0f, num_segments = 0, thickness = 1.0f
@[c:'ImDrawList_AddEllipseEx']
fn im_draw_list_add_ellipse_ex(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32, rot f32, num_segments int, thickness f32)

@[c:'ImDrawList_AddEllipseFilled']
fn im_draw_list_add_ellipse_filled(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32)

// Implied rot = 0.0f, num_segments = 0
@[c:'ImDrawList_AddEllipseFilledEx']
fn im_draw_list_add_ellipse_filled_ex(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32, rot f32, num_segments int)

@[c:'ImDrawList_AddText']
fn im_draw_list_add_text(self &ImDrawList, pos ImVec2, col ImU32, text_begin &i8)

// Implied text_end = NULL
@[c:'ImDrawList_AddTextEx']
fn im_draw_list_add_text_ex(self &ImDrawList, pos ImVec2, col ImU32, text_begin &i8, text_end &i8)

@[c:'ImDrawList_AddTextImFontPtr']
fn im_draw_list_add_text_im_font_ptr(self &ImDrawList, font &ImFont, font_size f32, pos ImVec2, col ImU32, text_begin &i8)

// Implied text_end = NULL, wrap_width = 0.0f, cpu_fine_clip_rect = NULL
@[c:'ImDrawList_AddTextImFontPtrEx']
fn im_draw_list_add_text_im_font_ptr_ex(self &ImDrawList, font &ImFont, font_size f32, pos ImVec2, col ImU32, text_begin &i8, text_end &i8, wrap_width f32, cpu_fine_clip_rect &C.ImVec4)

@[c:'ImDrawList_AddBezierCubic']
fn im_draw_list_add_bezier_cubic(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32, thickness f32, num_segments int)

// Cubic Bezier (4 control points)
@[c:'ImDrawList_AddBezierQuadratic']
fn im_draw_list_add_bezier_quadratic(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32, thickness f32, num_segments int)

// Quadratic Bezier (3 control points)
// General polygon
// - Only simple polygons are supported by filling functions (no self-intersections, no holes).
// - Concave polygon fill is more expensive than convex one: it has O(N^2) complexity. Provided as a convenience for the user but not used by the main library.
@[c:'ImDrawList_AddPolyline']
fn im_draw_list_add_polyline(self &ImDrawList, points &ImVec2, num_points int, col ImU32, flags ImDrawFlags, thickness f32)

@[c:'ImDrawList_AddConvexPolyFilled']
fn im_draw_list_add_convex_poly_filled(self &ImDrawList, points &ImVec2, num_points int, col ImU32)

@[c:'ImDrawList_AddConcavePolyFilled']
fn im_draw_list_add_concave_poly_filled(self &ImDrawList, points &ImVec2, num_points int, col ImU32)

// Image primitives
// - Read FAQ to understand what ImTextureID is.
// - "p_min" and "p_max" represent the upper-left and lower-right corners of the rectangle.
// - "uv_min" and "uv_max" represent the normalized texture coordinates to use for those corners. Using (0,0)->(1,1) texture coordinates will generally display the entire texture.
@[c:'ImDrawList_AddImage']
fn im_draw_list_add_image(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2)

// Implied uv_min = ImVec2(0, 0), uv_max = ImVec2(1, 1), col = IM_COL32_WHITE
@[c:'ImDrawList_AddImageEx']
fn im_draw_list_add_image_ex(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2, uv_min ImVec2, uv_max ImVec2, col ImU32)

@[c:'ImDrawList_AddImageQuad']
fn im_draw_list_add_image_quad(self &ImDrawList, user_texture_id ImTextureID, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2)

// Implied uv1 = ImVec2(0, 0), uv2 = ImVec2(1, 0), uv3 = ImVec2(1, 1), uv4 = ImVec2(0, 1), col = IM_COL32_WHITE
@[c:'ImDrawList_AddImageQuadEx']
fn im_draw_list_add_image_quad_ex(self &ImDrawList, user_texture_id ImTextureID, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, uv1 ImVec2, uv2 ImVec2, uv3 ImVec2, uv4 ImVec2, col ImU32)

@[c:'ImDrawList_AddImageRounded']
fn im_draw_list_add_image_rounded(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2, uv_min ImVec2, uv_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags)

// Stateful path API, add points then finish with PathFillConvex() or PathStroke()
// - Important: filled shapes must always use clockwise winding order! The anti-aliasing fringe depends on it. Counter-clockwise shapes will have "inward" anti-aliasing.
//   so e.g. 'PathArcTo(center, radius, PI * -0.5f, PI)' is ok, whereas 'PathArcTo(center, radius, PI, PI * -0.5f)' won't have correct anti-aliasing when followed by PathFillConvex().
@[c:'ImDrawList_PathClear']
fn im_draw_list_path_clear(self &ImDrawList)

@[c:'ImDrawList_PathLineTo']
fn im_draw_list_path_line_to(self &ImDrawList, pos ImVec2)

@[c:'ImDrawList_PathLineToMergeDuplicate']
fn im_draw_list_path_line_to_merge_duplicate(self &ImDrawList, pos ImVec2)

@[c:'ImDrawList_PathFillConvex']
fn im_draw_list_path_fill_convex(self &ImDrawList, col ImU32)

@[c:'ImDrawList_PathFillConcave']
fn im_draw_list_path_fill_concave(self &ImDrawList, col ImU32)

@[c:'ImDrawList_PathStroke']
fn im_draw_list_path_stroke(self &ImDrawList, col ImU32, flags ImDrawFlags, thickness f32)

@[c:'ImDrawList_PathArcTo']
fn im_draw_list_path_arc_to(self &ImDrawList, center ImVec2, radius f32, a_min f32, a_max f32, num_segments int)

@[c:'ImDrawList_PathArcToFast']
fn im_draw_list_path_arc_to_fast(self &ImDrawList, center ImVec2, radius f32, a_min_of_12 int, a_max_of_12 int)

// Use precomputed angles for a 12 steps circle
@[c:'ImDrawList_PathEllipticalArcTo']
fn im_draw_list_path_elliptical_arc_to(self &ImDrawList, center ImVec2, radius ImVec2, rot f32, a_min f32, a_max f32)

// Implied num_segments = 0
@[c:'ImDrawList_PathEllipticalArcToEx']
fn im_draw_list_path_elliptical_arc_to_ex(self &ImDrawList, center ImVec2, radius ImVec2, rot f32, a_min f32, a_max f32, num_segments int)

// Ellipse
@[c:'ImDrawList_PathBezierCubicCurveTo']
fn im_draw_list_path_bezier_cubic_curve_to(self &ImDrawList, p2 ImVec2, p3 ImVec2, p4 ImVec2, num_segments int)

// Cubic Bezier (4 control points)
@[c:'ImDrawList_PathBezierQuadraticCurveTo']
fn im_draw_list_path_bezier_quadratic_curve_to(self &ImDrawList, p2 ImVec2, p3 ImVec2, num_segments int)

// Quadratic Bezier (3 control points)
@[c:'ImDrawList_PathRect']
fn im_draw_list_path_rect(self &ImDrawList, rect_min ImVec2, rect_max ImVec2, rounding f32, flags ImDrawFlags)

// Advanced: Draw Callbacks
// - May be used to alter render state (change sampler, blending, current shader). May be used to emit custom rendering commands (difficult to do correctly, but possible).
// - Use special ImDrawCallback_ResetRenderState callback to instruct backend to reset its render state to the default.
// - Your rendering loop must check for 'UserCallback' in ImDrawCmd and call the function instead of rendering triangles. All standard backends are honoring this.
// - For some backends, the callback may access selected render-states exposed by the backend in a ImplXXXX_RenderState structure pointed to by platform_io.Renderer_RenderState.
// - IMPORTANT: please be mindful of the different level of indirection between using size==0 (copying argument) and using size>0 (copying pointed data into a buffer).
//   - If userdata_size == 0: we copy/store the 'userdata' argument as-is. It will be available unmodified in ImDrawCmd::UserCallbackData during render.
//   - If userdata_size > 0,  we copy/store 'userdata_size' bytes pointed to by 'userdata'. We store them in a buffer stored inside the drawlist. ImDrawCmd::UserCallbackData will point inside that buffer so you have to retrieve data from there. Your callback may need to use ImDrawCmd::UserCallbackDataSize if you expect dynamically-sized data.
//   - Support for userdata_size > 0 was added in v1.91.4, October 2024. So earlier code always only allowed to copy/store a simple void*.
@[c:'ImDrawList_AddCallback']
fn im_draw_list_add_callback(self &ImDrawList, callback ImDrawCallback, userdata voidptr)

// Implied userdata_size = 0
@[c:'ImDrawList_AddCallbackEx']
fn im_draw_list_add_callback_ex(self &ImDrawList, callback ImDrawCallback, userdata voidptr, userdata_size usize)

// Advanced: Miscellaneous
@[c:'ImDrawList_AddDrawCmd']
fn im_draw_list_add_draw_cmd(self &ImDrawList)

// This is useful if you need to forcefully create a new draw call (to allow for dependent rendering / blending). Otherwise primitives are merged into the same draw-call as much as possible
@[c:'ImDrawList_CloneOutput']
fn im_draw_list_clone_output(self &ImDrawList) &ImDrawList

// Create a clone of the CmdBuffer/IdxBuffer/VtxBuffer.
// Advanced: Channels
// - Use to split render into layers. By switching channels to can render out-of-order (e.g. submit FG primitives before BG primitives)
// - Use to minimize draw calls (e.g. if going back-and-forth between multiple clipping rectangles, prefer to append into separate channels then merge at the end)
// - This API shouldn't have been in ImDrawList in the first place!
//   Prefer using your own persistent instance of ImDrawListSplitter as you can stack them.
//   Using the ImDrawList::ChannelsXXXX you cannot stack a split over another.
@[c:'ImDrawList_ChannelsSplit']
fn im_draw_list_channels_split(self &ImDrawList, count int)

@[c:'ImDrawList_ChannelsMerge']
fn im_draw_list_channels_merge(self &ImDrawList)

@[c:'ImDrawList_ChannelsSetCurrent']
fn im_draw_list_channels_set_current(self &ImDrawList, n int)

// Advanced: Primitives allocations
// - We render triangles (three vertices)
// - All primitives needs to be reserved via PrimReserve() beforehand.
@[c:'ImDrawList_PrimReserve']
fn im_draw_list_prim_reserve(self &ImDrawList, idx_count int, vtx_count int)

@[c:'ImDrawList_PrimUnreserve']
fn im_draw_list_prim_unreserve(self &ImDrawList, idx_count int, vtx_count int)

@[c:'ImDrawList_PrimRect']
fn im_draw_list_prim_rect(self &ImDrawList, a ImVec2, b ImVec2, col ImU32)

// Axis aligned rectangle (composed of two triangles)
@[c:'ImDrawList_PrimRectUV']
fn im_draw_list_prim_rect_uv(self &ImDrawList, a ImVec2, b ImVec2, uv_a ImVec2, uv_b ImVec2, col ImU32)

@[c:'ImDrawList_PrimQuadUV']
fn im_draw_list_prim_quad_uv(self &ImDrawList, a ImVec2, b ImVec2, c ImVec2, d ImVec2, uv_a ImVec2, uv_b ImVec2, uv_c ImVec2, uv_d ImVec2, col ImU32)

@[c:'ImDrawList_PrimWriteVtx']
fn im_draw_list_prim_write_vtx(self &ImDrawList, pos ImVec2, uv ImVec2, col ImU32)

@[c:'ImDrawList_PrimWriteIdx']
fn im_draw_list_prim_write_idx(self &ImDrawList, idx ImDrawIdx)

@[c:'ImDrawList_PrimVtx']
fn im_draw_list_prim_vtx(self &ImDrawList, pos ImVec2, uv ImVec2, col ImU32)

// Write vertex with unique index
// [Internal helpers]
@[c:'ImDrawList__ResetForNewFrame']
fn im_draw_list__reset_for_new_frame(self &ImDrawList)

@[c:'ImDrawList__ClearFreeMemory']
fn im_draw_list__clear_free_memory(self &ImDrawList)

@[c:'ImDrawList__PopUnusedDrawCmd']
fn im_draw_list__pop_unused_draw_cmd(self &ImDrawList)

@[c:'ImDrawList__TryMergeDrawCmds']
fn im_draw_list__try_merge_draw_cmds(self &ImDrawList)

@[c:'ImDrawList__OnChangedClipRect']
fn im_draw_list__on_changed_clip_rect(self &ImDrawList)

@[c:'ImDrawList__OnChangedTextureID']
fn im_draw_list__on_changed_texture_id(self &ImDrawList)

@[c:'ImDrawList__OnChangedVtxOffset']
fn im_draw_list__on_changed_vtx_offset(self &ImDrawList)

@[c:'ImDrawList__SetTextureID']
fn im_draw_list__set_texture_id(self &ImDrawList, texture_id ImTextureID)

@[c:'ImDrawList__CalcCircleAutoSegmentCount']
fn im_draw_list__calc_circle_auto_segment_count(self &ImDrawList, radius f32) int

@[c:'ImDrawList__PathArcToFastEx']
fn im_draw_list__path_arc_to_fast_ex(self &ImDrawList, center ImVec2, radius f32, a_min_sample int, a_max_sample int, a_step int)

@[c:'ImDrawList__PathArcToN']
fn im_draw_list__path_arc_to_n(self &ImDrawList, center ImVec2, radius f32, a_min f32, a_max f32, num_segments int)

// All draw data to render a Dear ImGui frame
// (NB: the style and the naming convention here is a little inconsistent, we currently preserve them for backward compatibility purpose,
// as this is one of the oldest structure exposed by the library! Basically, ImDrawList == CmdList)
struct ImDrawData { 
	valid bool
// Only valid after Render() is called and before the next NewFrame() is called.
	cmdListsCount int
// Number of ImDrawList* to render (should always be == CmdLists.size)
	totalIdxCount int
// For convenience, sum of all ImDrawList's IdxBuffer.Size
	totalVtxCount int
// For convenience, sum of all ImDrawList's VtxBuffer.Size
	cmdLists ImVector_ImDrawListPtr
// Array of ImDrawList* to render. The ImDrawLists are owned by C.ImGuiContext and only pointed to from here.
	displayPos ImVec2
// Top-left position of the viewport to render (== top-left of the orthogonal projection matrix to use) (== GetMainViewport()->Pos for the main viewport, == (0.0) in most single-viewport applications)
	displaySize ImVec2
// Size of the viewport to render (== GetMainViewport()->Size for the main viewport, == io.DisplaySize in most single-viewport applications)
	framebufferScale ImVec2
// Amount of pixels for each unit of DisplaySize. Based on io.DisplayFramebufferScale. Generally (1,1) on normal display, (2,2) on OSX with Retina display.
	ownerViewport &ImGuiViewport
}
@[c:'ImDrawData_Clear']
fn im_draw_data_clear(self &ImDrawData)

@[c:'ImDrawData_AddDrawList']
fn im_draw_data_add_draw_list(self &ImDrawData, draw_list &ImDrawList)

// Helper to add an external draw list into an existing ImDrawData.
@[c:'ImDrawData_DeIndexAllBuffers']
fn im_draw_data_de_index_all_buffers(self &ImDrawData)

// Helper to convert all buffers from indexed to non-indexed, in case you cannot render indexed. Note: this is slow and most likely a waste of resources. Always prefer indexed rendering!
@[c:'ImDrawData_ScaleClipRects']
fn im_draw_data_scale_clip_rects(self &ImDrawData, fb_scale ImVec2)

// Helper to scale the ClipRect field of each ImDrawCmd. Use if your final output buffer is at a different scale than Dear ImGui expects, or if there is a difference between your window resolution and framebuffer resolution.
//-----------------------------------------------------------------------------
// [SECTION] Font API (ImFontConfig, ImFontGlyph, ImFontAtlasFlags, ImFontAtlas, ImFontGlyphRangesBuilder, ImFont)
//-----------------------------------------------------------------------------
// A font input/source (we may rename this to ImFontSource in the future)
struct ImFontConfig { 
	fontData voidptr
//          // TTF/OTF data
	fontDataSize int
//          // TTF/OTF data size
	fontDataOwnedByAtlas bool
// true     // TTF/OTF data ownership taken by the container ImFontAtlas (will delete memory itself).
	mergeMode bool
// false    // Merge into previous ImFont, so you can combine multiple inputs font into one ImFont (e.g. ASCII font + icons + Japanese glyphs). You may want to use GlyphOffset.y when merge font of different heights.
	pixelSnapH bool
// false    // Align every glyph AdvanceX to pixel boundaries. Useful e.g. if you are merging a non-pixel aligned font with the default font. If enabled, you can set OversampleH/V to 1.
	fontNo int
// 0        // Index of font within TTF/OTF file
	oversampleH int
// 0 (2)    // Rasterize at higher quality for sub-pixel positioning. 0 == auto == 1 or 2 depending on size. Note the difference between 2 and 3 is minimal. You can reduce this to 1 for large glyphs save memory. Read https://github.com/nothings/stb/blob/master/tests/oversample/README.md for details.
	oversampleV int
// 0 (1)    // Rasterize at higher quality for sub-pixel positioning. 0 == auto == 1. This is not really useful as we don't use sub-pixel positions on the Y axis.
	sizePixels f32
//          // Size in pixels for rasterizer (more or less maps to the resulting font height).
//ImVec2        GlyphExtraSpacing;      // 0, 0     // (REMOVED IN 1.91.9: use GlyphExtraAdvanceX)
	glyphOffset ImVec2
// 0, 0     // Offset all glyphs from this font input.
	glyphRanges &C.ImWchar
// NULL     // THE ARRAY DATA NEEDS TO PERSIST AS LONG AS THE FONT IS ALIVE. Pointer to a user-provided list of Unicode range (2 value per range, values are inclusive, zero-terminated list).
	glyphMinAdvanceX f32
// 0        // Minimum AdvanceX for glyphs, set Min to align font icons, set both Min/Max to enforce mono-space font
	glyphMaxAdvanceX f32
// FLT_MAX  // Maximum AdvanceX for glyphs
	glyphExtraAdvanceX f32
// 0        // Extra spacing (in pixels) between glyphs. Please contact us if you are using this.
	fontBuilderFlags u32
// 0        // Settings for custom font builder. THIS IS BUILDER IMPLEMENTATION DEPENDENT. Leave as zero if unsure.
	rasterizerMultiply f32
// 1.0f     // Linearly brighten (>1.0f) or darken (<1.0f) font output. Brightening small fonts may be a good workaround to make them more readable. This is a silly thing we may remove in the future.
	rasterizerDensity f32
// 1.0f     // DPI scale for rasterization, not altering other font metrics: make it easy to swap between e.g. a 100% and a 400% fonts for a zooming display. IMPORTANT: If you increase this it is expected that you increase font scale accordingly, otherwise quality may look lowered.
	ellipsisChar C.ImWchar
// 0        // Explicitly specify Unicode codepoint of ellipsis character. When fonts are being merged first specified ellipsis will be used.
// [Internal]
	name [40]i8
// Name (strictly to ease debugging)
	dstFont &ImFont
}
// Hold rendering data for one glyph.
// (Note: some language parsers may fail to convert the 31+1 bitfield members, in this case maybe drop store a single u32 or we can rework this)
struct ImFontGlyph { 
	colored u32
// Flag to indicate glyph is colored and should generally ignore tinting (make it usable with no shift on little-endian as this is used in loops)
	visible u32
// Flag to indicate glyph has no visible pixels (e.g. space). Allow early out when rendering.
	codepoint u32
// 0x0000..0x10FFFF
	advanceX f32
// Horizontal distance to advance layout with
	x0 f32
	y0 f32
	x1 f32
	y1 f32
// Glyph corners
	u0 f32
	v0 f32
	u1 f32
	v1 f32
}
// Helper to build glyph ranges from text/string data. Feed your application strings/characters to it then call BuildRanges().
// This is essentially a tightly packed of vector of 64k booleans = 8KB storage.
struct ImFontGlyphRangesBuilder { 
	usedChars ImVector_ImU32
}
@[c:'ImFontGlyphRangesBuilder_Clear']
fn im_font_glyph_ranges_builder_clear(self &ImFontGlyphRangesBuilder)

@[c:'ImFontGlyphRangesBuilder_GetBit']
fn im_font_glyph_ranges_builder_get_bit(self &ImFontGlyphRangesBuilder, n usize) bool

// Get bit n in the array
@[c:'ImFontGlyphRangesBuilder_SetBit']
fn im_font_glyph_ranges_builder_set_bit(self &ImFontGlyphRangesBuilder, n usize)

// Set bit n in the array
@[c:'ImFontGlyphRangesBuilder_AddChar']
fn im_font_glyph_ranges_builder_add_char(self &ImFontGlyphRangesBuilder, c C.ImWchar)

// Add character
@[c:'ImFontGlyphRangesBuilder_AddText']
fn im_font_glyph_ranges_builder_add_text(self &ImFontGlyphRangesBuilder, text &i8, text_end &i8)

// Add string (each character of the UTF-8 string are added)
@[c:'ImFontGlyphRangesBuilder_AddRanges']
fn im_font_glyph_ranges_builder_add_ranges(self &ImFontGlyphRangesBuilder, ranges &C.ImWchar)

// Add ranges, e.g. builder.AddRanges(ImFontAtlas::GetGlyphRangesDefault()) to force add all of ASCII/Latin+Ext
@[c:'ImFontGlyphRangesBuilder_BuildRanges']
fn im_font_glyph_ranges_builder_build_ranges(self &ImFontGlyphRangesBuilder, out_ranges &ImVector_ImWchar)

// Output new ranges (ImVector_Construct()/ImVector_Destruct() can be used to safely construct out_ranges)
// See ImFontAtlas::AddCustomRectXXX functions.
struct ImFontAtlasCustomRect { 
	x u16
	y u16
// Output   // Packed position in Atlas
// [Internal]
	width u16
	height u16
// Input    // Desired rectangle dimension
	glyphID u32
// Input    // For custom font glyphs only (ID < 0x110000)
	glyphColored u32
// Input  // For custom font glyphs only: glyph is colored, removed tinting.
	glyphAdvanceX f32
// Input    // For custom font glyphs only: glyph xadvance
	glyphOffset ImVec2
// Input    // For custom font glyphs only: glyph display offset
	font &ImFont
}
@[c:'ImFontAtlasCustomRect_IsPacked']
fn im_font_atlas_custom_rect_is_packed(self &ImFontAtlasCustomRect) bool

// Flags for ImFontAtlas build
enum ImFontAtlasFlags_ {
	none = 0
	no_power_of_two_height = 1 << 0
// Don't round the height to next power of two
	no_mouse_cursors = 1 << 1
// Don't build software mouse cursors into the atlas (save a little texture memory)
	no_baked_lines = 1 << 2
}

// Load and rasterize multiple TTF/OTF fonts into a same texture. The font atlas will build a single texture holding:
//  - One or more fonts.
//  - Custom graphics data needed to render the shapes needed by Dear ImGui.
//  - Mouse cursor shapes for software cursor rendering (unless setting 'Flags |= ImFontAtlasFlags_NoMouseCursors' in the font atlas).
// It is the user-code responsibility to setup/build the atlas, then upload the pixel data into a texture accessible by your graphics api.
//  - Optionally, call any of the AddFont*** functions. If you don't call any, the default font embedded in the code will be loaded for you.
//  - Call GetTexDataAsAlpha8() or GetTexDataAsRGBA32() to build and retrieve pixels data.
//  - Upload the pixels data into a texture within your graphics system (see imgui_impl_xxxx.cpp examples)
//  - Call SetTexID(my_tex_id); and pass the pointer/identifier to your texture in a format natural to your graphics API.
//    This value will be passed back to you during rendering to identify the texture. Read FAQ entry about ImTextureID for more details.
// Common pitfalls:
// - If you pass a 'glyph_ranges' array to AddFont*** functions, you need to make sure that your array persist up until the
//   atlas is build (when calling GetTexData*** or Build()). We only copy the pointer, not the data.
// - Important: By default, AddFontFromMemoryTTF() takes ownership of the data. Even though we are not writing to it, we will free the pointer on destruction.
//   You can set font_cfg->FontDataOwnedByAtlas=false to keep ownership of your data and it won't be freed,
// - Even though many functions are suffixed with "TTF", OTF data is supported just as well.
// - This is an old API and it is currently awkward for those and various other reasons! We will address them in the future!
struct ImFontAtlas { 
//-------------------------------------------
// Glyph Ranges
//-------------------------------------------
//-------------------------------------------
// [ALPHA] Custom Rectangles/Glyphs API
//-------------------------------------------
//-------------------------------------------
// Members
//-------------------------------------------
// Input
	flags ImFontAtlasFlags
// Build flags (see ImFontAtlasFlags_)
	texID ImTextureID
// User data to refer to the texture once it has been uploaded to user's graphic systems. It is passed back to you during rendering via the ImDrawCmd structure.
	texDesiredWidth int
// Texture width desired by user before Build(). Must be a power-of-two. If have many glyphs your graphics API have texture size restrictions you may want to increase texture width to decrease height.
	texGlyphPadding int
// FIXME: Should be called "TexPackPadding". Padding between glyphs within texture in pixels. Defaults to 1. If your rendering method doesn't rely on bilinear filtering you may set this to 0 (will also need to set AntiAliasedLinesUseTex = false).
	userData voidptr
// Store your own atlas related user-data (if e.g. you have multiple font atlas).
// [Internal]
// NB: Access texture data via GetTexData*() calls! Which will setup a default font for you.
	locked bool
// Marked as Locked by ImGui::NewFrame() so attempt to modify the atlas will assert.
	texReady bool
// Set when texture was built matching current font input
	texPixelsUseColors bool
// Tell whether our texture data is known to use colors (rather than just alpha channel), in order to help backend select a format.
	texPixelsAlpha8 &u8
// 1 component per pixel, each component is unsigned 8-bit. Total size = TexWidth * TexHeight
	texPixelsRGBA32 &u32
// 4 component per pixel, each component is unsigned 8-bit. Total size = TexWidth * TexHeight * 4
	texWidth int
// Texture width calculated during Build().
	texHeight int
// Texture height calculated during Build().
	texUvScale ImVec2
// = (1.0f/TexWidth, 1.0f/TexHeight)
	texUvWhitePixel ImVec2
// Texture coordinates to a white pixel
	fonts ImVector_ImFontPtr
// Hold all the fonts returned by AddFont*. Fonts[0] is the default font upon calling ImGui::NewFrame(), use ImGui::PushFont()/PopFont() to change the current font.
	customRects ImVector_ImFontAtlasCustomRect
// Rectangles for packing custom texture data into the atlas.
	sources ImVector_ImFontConfig
// Source/configuration data
	texUvLines [33]C.ImVec4
// UVs for baked anti-aliased lines
// [Internal] Font builder
	fontBuilderIO &C.ImFontBuilderIO
// Opaque interface to a font builder (default to stb_truetype, can be changed to use FreeType by defining IMGUI_ENABLE_FREETYPE).
	fontBuilderFlags u32
// Shared flags (for all fonts) for custom font builder. THIS IS BUILD IMPLEMENTATION DEPENDENT. Per-font override is also available in ImFontConfig.
// [Internal] Packing data
	packIdMouseCursors int
// Custom texture rectangle ID for white pixel and mouse cursors
	packIdLines int
// Custom texture rectangle ID for baked anti-aliased lines
// [Obsolete]
//typedef ImFontAtlasCustomRect    CustomRect;              // OBSOLETED in 1.72+
}
@[c:'ImFontAtlas_AddFont']
fn im_font_atlas_add_font(self &ImFontAtlas, font_cfg &ImFontConfig) &ImFont

@[c:'ImFontAtlas_AddFontDefault']
fn im_font_atlas_add_font_default(self &ImFontAtlas, font_cfg &ImFontConfig) &ImFont

@[c:'ImFontAtlas_AddFontFromFileTTF']
fn im_font_atlas_add_font_from_file_ttf(self &ImFontAtlas, filename &i8, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

@[c:'ImFontAtlas_AddFontFromMemoryTTF']
fn im_font_atlas_add_font_from_memory_ttf(self &ImFontAtlas, font_data voidptr, font_data_size int, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

// Note: Transfer ownership of 'ttf_data' to ImFontAtlas! Will be deleted after destruction of the atlas. Set font_cfg->FontDataOwnedByAtlas=false to keep ownership of your data and it won't be freed.
@[c:'ImFontAtlas_AddFontFromMemoryCompressedTTF']
fn im_font_atlas_add_font_from_memory_compressed_ttf(self &ImFontAtlas, compressed_font_data voidptr, compressed_font_data_size int, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

// 'compressed_font_data' still owned by caller. Compress with binary_to_compressed_c.cpp.
@[c:'ImFontAtlas_AddFontFromMemoryCompressedBase85TTF']
fn im_font_atlas_add_font_from_memory_compressed_base85_ttf(self &ImFontAtlas, compressed_font_data_base85 &i8, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &C.ImWchar) &ImFont

// 'compressed_font_data_base85' still owned by caller. Compress with binary_to_compressed_c.cpp with -base85 parameter.
@[c:'ImFontAtlas_ClearInputData']
fn im_font_atlas_clear_input_data(self &ImFontAtlas)

// Clear input data (all ImFontConfig structures including sizes, TTF data, glyph ranges, etc.) = all the data used to build the texture and fonts.
@[c:'ImFontAtlas_ClearFonts']
fn im_font_atlas_clear_fonts(self &ImFontAtlas)

// Clear input+output font data (same as ClearInputData() + glyphs storage, UV coordinates).
@[c:'ImFontAtlas_ClearTexData']
fn im_font_atlas_clear_tex_data(self &ImFontAtlas)

// Clear output texture data (CPU side). Saves RAM once the texture has been copied to graphics memory.
@[c:'ImFontAtlas_Clear']
fn im_font_atlas_clear(self &ImFontAtlas)

// Clear all input and output.
// Build atlas, retrieve pixel data.
// User is in charge of copying the pixels into graphics memory (e.g. create a texture with your engine). Then store your texture handle with SetTexID().
// The pitch is always = Width * BytesPerPixels (1 or 4)
// Building in RGBA32 format is provided for convenience and compatibility, but note that unless you manually manipulate or copy color data into
// the texture (e.g. when using the AddCustomRect*** api), then the RGB pixels emitted will always be white (~75% of memory/bandwidth waste.
@[c:'ImFontAtlas_Build']
fn im_font_atlas_build(self &ImFontAtlas) bool

// Build pixels data. This is called automatically for you by the GetTexData*** functions.
@[c:'ImFontAtlas_GetTexDataAsAlpha8']
fn im_font_atlas_get_tex_data_as_alpha8(self &ImFontAtlas, out_pixels &&u8, out_width &int, out_height &int, out_bytes_per_pixel &int)

// 1 byte per-pixel
@[c:'ImFontAtlas_GetTexDataAsRGBA32']
fn im_font_atlas_get_tex_data_as_rgba_32(self &ImFontAtlas, out_pixels &&u8, out_width &int, out_height &int, out_bytes_per_pixel &int)

// 4 bytes-per-pixel
@[c:'ImFontAtlas_IsBuilt']
fn im_font_atlas_is_built(self &ImFontAtlas) bool

// Bit ambiguous: used to detect when user didn't build texture but effectively we should check TexID != 0 except that would be backend dependent...
@[c:'ImFontAtlas_SetTexID']
fn im_font_atlas_set_tex_id(self &ImFontAtlas, id ImTextureID)

// Helpers to retrieve list of common Unicode ranges (2 value per range, values are inclusive, zero-terminated list)
// NB: Make sure that your string are UTF-8 and NOT in your local code page.
// Read https://github.com/ocornut/imgui/blob/master/docs/FONTS.md/#about-utf-8-encoding for details.
// NB: Consider using ImFontGlyphRangesBuilder to build glyph ranges from textual data.
@[c:'ImFontAtlas_GetGlyphRangesDefault']
fn im_font_atlas_get_glyph_ranges_default(self &ImFontAtlas) &C.ImWchar

// Basic Latin, Extended Latin
@[c:'ImFontAtlas_GetGlyphRangesGreek']
fn im_font_atlas_get_glyph_ranges_greek(self &ImFontAtlas) &C.ImWchar

// Default + Greek and Coptic
@[c:'ImFontAtlas_GetGlyphRangesKorean']
fn im_font_atlas_get_glyph_ranges_korean(self &ImFontAtlas) &C.ImWchar

// Default + Korean characters
@[c:'ImFontAtlas_GetGlyphRangesJapanese']
fn im_font_atlas_get_glyph_ranges_japanese(self &ImFontAtlas) &C.ImWchar

// Default + Hiragana, Katakana, Half-Width, Selection of 2999 Ideographs
@[c:'ImFontAtlas_GetGlyphRangesChineseFull']
fn im_font_atlas_get_glyph_ranges_chinese_full(self &ImFontAtlas) &C.ImWchar

// Default + Half-Width + Japanese Hiragana/Katakana + full set of about 21000 CJK Unified Ideographs
@[c:'ImFontAtlas_GetGlyphRangesChineseSimplifiedCommon']
fn im_font_atlas_get_glyph_ranges_chinese_simplified_common(self &ImFontAtlas) &C.ImWchar

// Default + Half-Width + Japanese Hiragana/Katakana + set of 2500 CJK Unified Ideographs for common simplified Chinese
@[c:'ImFontAtlas_GetGlyphRangesCyrillic']
fn im_font_atlas_get_glyph_ranges_cyrillic(self &ImFontAtlas) &C.ImWchar

// Default + about 400 Cyrillic characters
@[c:'ImFontAtlas_GetGlyphRangesThai']
fn im_font_atlas_get_glyph_ranges_thai(self &ImFontAtlas) &C.ImWchar

// Default + Thai characters
@[c:'ImFontAtlas_GetGlyphRangesVietnamese']
fn im_font_atlas_get_glyph_ranges_vietnamese(self &ImFontAtlas) &C.ImWchar

// Default + Vietnamese characters
// You can request arbitrary rectangles to be packed into the atlas, for your own purposes.
// - After calling Build(), you can query the rectangle position and render your pixels.
// - If you render colored output, set 'atlas->TexPixelsUseColors = true' as this may help some backends decide of preferred texture format.
// - You can also request your rectangles to be mapped as font glyph (given a font + Unicode point),
//   so you can render e.g. custom colorful icons and use them as regular glyphs.
// - Read docs/FONTS.md for more details about using colorful icons.
// - Note: this API may be redesigned later in order to support multi-monitor varying DPI settings.
@[c:'ImFontAtlas_AddCustomRectRegular']
fn im_font_atlas_add_custom_rect_regular(self &ImFontAtlas, width int, height int) int

@[c:'ImFontAtlas_AddCustomRectFontGlyph']
fn im_font_atlas_add_custom_rect_font_glyph(self &ImFontAtlas, font &ImFont, id C.ImWchar, width int, height int, advance_x f32, offset ImVec2) int

@[c:'ImFontAtlas_GetCustomRectByIndex']
fn im_font_atlas_get_custom_rect_by_index(self &ImFontAtlas, index int) &ImFontAtlasCustomRect

// [Internal]
@[c:'ImFontAtlas_CalcCustomRectUV']
fn im_font_atlas_calc_custom_rect_uv(self &ImFontAtlas, rect &ImFontAtlasCustomRect, out_uv_min &ImVec2, out_uv_max &ImVec2)

// Font runtime data and rendering
// ImFontAtlas automatically loads a default embedded font for you when you call GetTexDataAsAlpha8() or GetTexDataAsRGBA32().
struct ImFont { 
// [Internal] Members: Hot ~20/24 bytes (for CalcTextSize)
	indexAdvanceX ImVector_float
// 12-16 // out // Sparse. Glyphs->AdvanceX in a directly indexable way (cache-friendly for CalcTextSize functions which only this info, and are often bottleneck in large UI).
	fallbackAdvanceX f32
// 4     // out // = FallbackGlyph->AdvanceX
	fontSize f32
// 4     // in  // Height of characters/line, set during loading (don't change after loading)
// [Internal] Members: Hot ~28/40 bytes (for RenderText loop)
	indexLookup ImVector_ImU16
// 12-16 // out // Sparse. Index glyphs by Unicode code-point.
	glyphs ImVector_ImFontGlyph
// 12-16 // out // All glyphs.
	fallbackGlyph &ImFontGlyph
// 4-8   // out // = FindGlyph(FontFallbackChar)
// [Internal] Members: Cold ~32/40 bytes
// Conceptually Sources[] is the list of font sources merged to create this font.
	containerAtlas &ImFontAtlas
// 4-8   // out // What we has been loaded into
	sources &ImFontConfig
// 4-8   // in  // Pointer within ContainerAtlas->Sources[], to SourcesCount instances
	sourcesCount i16
// 2     // in  // Number of ImFontConfig involved in creating this font. Usually 1, or >1 when merging multiple font sources into one ImFont.
	ellipsisCharCount i16
// 1     // out // 1 or 3
	ellipsisChar C.ImWchar
// 2-4   // out // Character used for ellipsis rendering ('...').
	fallbackChar C.ImWchar
// 2-4   // out // Character used if a glyph isn't found (U+FFFD, '?')
	ellipsisWidth f32
// 4     // out // Total ellipsis Width
	ellipsisCharStep f32
// 4     // out // Step between characters when EllipsisCount > 0
	scale f32
// 4     // in  // Base font scale (1.0f), multiplied by the per-window font scale which you can adjust with SetWindowFontScale()
	ascent f32
	descent f32
// 4+4   // out // Ascent: distance from top to bottom of e.g. 'A' [0..FontSize] (unscaled)
	metricsTotalSurface int
// 4     // out // Total surface in pixels to get an idea of the font rasterization/texture cost (not exact, we approximate the cost of padding between glyphs)
	dirtyLookupTables bool
// 1     // out //
	used8kPagesMap [1]ImU8
}
@[c:'ImFont_FindGlyph']
fn im_font_find_glyph(self &ImFont, c C.ImWchar) &ImFontGlyph

@[c:'ImFont_FindGlyphNoFallback']
fn im_font_find_glyph_no_fallback(self &ImFont, c C.ImWchar) &ImFontGlyph

@[c:'ImFont_GetCharAdvance']
fn im_font_get_char_advance(self &ImFont, c C.ImWchar) f32

@[c:'ImFont_IsLoaded']
fn im_font_is_loaded(self &ImFont) bool

@[c:'ImFont_GetDebugName']
fn im_font_get_debug_name(self &ImFont) &i8

// [Internal] Don't use!
// 'max_width' stops rendering after a certain width (could be turned into a 2d size). FLT_MAX to disable.
// 'wrap_width' enable automatic word-wrapping across multiple lines to fit into given width. 0.0f to disable.
@[c:'ImFont_CalcTextSizeA']
fn im_font_calc_text_size_a(self &ImFont, size f32, max_width f32, wrap_width f32, text_begin &i8) ImVec2

// Implied text_end = NULL, remaining = NULL
@[c:'ImFont_CalcTextSizeAEx']
fn im_font_calc_text_size_ae_x(self &ImFont, size f32, max_width f32, wrap_width f32, text_begin &i8, text_end &i8, remaining &&u8) ImVec2

// utf8
@[c:'ImFont_CalcWordWrapPositionA']
fn im_font_calc_word_wrap_position_a(self &ImFont, scale f32, text &i8, text_end &i8, wrap_width f32) &i8

@[c:'ImFont_RenderChar']
fn im_font_render_char(self &ImFont, draw_list &ImDrawList, size f32, pos ImVec2, col ImU32, c C.ImWchar)

@[c:'ImFont_RenderText']
fn im_font_render_text(self &ImFont, draw_list &ImDrawList, size f32, pos ImVec2, col ImU32, clip_rect C.ImVec4, text_begin &i8, text_end &i8, wrap_width f32, cpu_fine_clip bool)

// [Internal] Don't use!
@[c:'ImFont_BuildLookupTable']
fn im_font_build_lookup_table(self &ImFont)

@[c:'ImFont_ClearOutputData']
fn im_font_clear_output_data(self &ImFont)

@[c:'ImFont_GrowIndex']
fn im_font_grow_index(self &ImFont, new_size int)

@[c:'ImFont_AddGlyph']
fn im_font_add_glyph(self &ImFont, src_cfg &ImFontConfig, c C.ImWchar, x0 f32, y0 f32, x1 f32, y1 f32, u0 f32, v0 f32, u1 f32, v1 f32, advance_x f32)

@[c:'ImFont_AddRemapChar']
fn im_font_add_remap_char(self &ImFont, dst C.ImWchar, src C.ImWchar, overwrite_dst bool)

// Makes 'dst' character/glyph points to 'src' character/glyph. Currently needs to be called AFTER fonts have been built.
@[c:'ImFont_IsGlyphRangeUnused']
fn im_font_is_glyph_range_unused(self &ImFont, c_begin u32, c_last u32) bool

//-----------------------------------------------------------------------------
// [SECTION] Viewports
//-----------------------------------------------------------------------------
// Flags stored in ImGuiViewport::Flags, giving indications to the platform backends.
enum ImGuiViewportFlags_ {
 viewport_flags_none = 0
 viewport_flags_is_platform_window = 1 << 0
// Represent a Platform Window
 viewport_flags_is_platform_monitor = 1 << 1
// Represent a Platform Monitor (unused yet)
 viewport_flags_owned_by_app = 1 << 2
}

// - Currently represents the Platform Window created by the application which is hosting our Dear ImGui windows.
// - In 'docking' branch with multi-viewport enabled, we extend this concept to have multiple active viewports.
// - In the future we will extend this concept further to also represent Platform Monitor and support a "no main platform window" operation mode.
// - About Main Area vs Work Area:
//   - Main Area = entire viewport.
//   - Work Area = entire viewport minus sections used by main menu bars (for platform windows), or by task bar (for platform monitor).
//   - Windows are generally trying to stay within the Work Area of their host viewport.
struct ImGuiViewport { 
	iD ID
// Unique identifier for the viewport
	flags ImGuiViewportFlags
// See ImGuiViewportFlags_
	pos ImVec2
// Main Area: Position of the viewport (Dear ImGui coordinates are the same as OS desktop/native coordinates)
	size ImVec2
// Main Area: Size of the viewport.
	workPos ImVec2
// Work Area: Position of the viewport minus task bars, menus bars, status bars (>= Pos)
	workSize ImVec2
// Work Area: Size of the viewport minus task bars, menu bars, status bars (<= Size)
// Platform/Backend Dependent Data
	platformHandle voidptr
// void* to hold higher-level, platform window handle (e.g. HWND, GLFWWindow*, SDL_Window*)
	platformHandleRaw voidptr
}
// Helpers
@[c:'ImGuiViewport_GetCenter']
fn viewport_get_center(self &ImGuiViewport) ImVec2

@[c:'ImGuiViewport_GetWorkCenter']
fn viewport_get_work_center(self &ImGuiViewport) ImVec2

//-----------------------------------------------------------------------------
// [SECTION] Platform Dependent Interfaces
//-----------------------------------------------------------------------------
// Access via ImGui::GetPlatformIO()
struct ImGuiPlatformIO { 
//------------------------------------------------------------------
// Input - Interface with OS and Platform backend (most common stuff)
//------------------------------------------------------------------
// Optional: Access OS clipboard
// (default to use native Win32 clipboard on Windows, otherwise uses a private clipboard. Override to access OS clipboard on other architectures)
	platform_GetClipboardTextFn fn (&C.ImGuiContext) &i8
	platform_SetClipboardTextFn fn (&C.ImGuiContext, &i8)
	platform_ClipboardUserData voidptr
// Optional: Open link/folder/file in OS Shell
// (default to use ShellExecuteW() on Windows, system() on Linux/Mac)
	platform_OpenInShellFn fn (&C.ImGuiContext, &i8) bool
	platform_OpenInShellUserData voidptr
// Optional: Notify OS Input Method Editor of the screen position of your cursor for text input position (e.g. when using Japanese/Chinese IME on Windows)
// (default to use native imm32 api on Windows)
	platform_SetImeDataFn fn (&C.ImGuiContext, &ImGuiViewport,  PlatformImeData)
	platform_ImeUserData voidptr
//void      (*SetPlatformImeDataFn)(ImGuiViewport* viewport, PlatformImeData* data); // [Renamed to platform_io.PlatformSetImeDataFn in 1.91.1]
// Optional: Platform locale
// [Experimental] Configure decimal point e.g. '.' or ',' useful for some languages (e.g. German), generally pulled from *localeconv()->decimal_point
	platform_LocaleDecimalPoint C.ImWchar
// '.'
//------------------------------------------------------------------
// Input - Interface with Renderer Backend
//------------------------------------------------------------------
// Written by some backends during ImplXXXX_RenderDrawData() call to point backend_specific ImplXXXX_RenderState* structure.
	renderer_RenderState voidptr
}
// (Optional) Support for IME (Input Method Editor) via the platform_io.Platform_SetImeDataFn() function.
struct PlatformImeData { 
	wantVisible bool
// A widget wants the IME to be visible
	inputPos ImVec2
// Position of the input cursor
	inputLineHeight f32
}
//-----------------------------------------------------------------------------
// [SECTION] Obsolete functions and types
// (Will be removed! Read 'API BREAKING CHANGES' section in imgui.cpp for details)
// Please keep your copy of dear imgui up to date! Occasionally set '#define IMGUI_DISABLE_OBSOLETE_FUNCTIONS' in imconfig.h to stay ahead.
//-----------------------------------------------------------------------------
// OBSOLETED in 1.91.9 (from February 2025)
@[c:'ImGui_ImageImVec4']
fn image_im_vec4(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, tint_col C.ImVec4, border_col C.ImVec4)

// <-- border_col was removed in favor of Col_ImageBorder.
// OBSOLETED in 1.91.0 (from July 2024)
@[c:'ImGui_PushButtonRepeat']
fn push_button_repeat(repeat bool)

@[c:'ImGui_PopButtonRepeat']
fn pop_button_repeat()

@[c:'ImGui_PushTabStop']
fn push_tab_stop(tab_stop bool)

@[c:'ImGui_PopTabStop']
fn pop_tab_stop()

@[c:'ImGui_GetContentRegionMax']
fn get_content_region_max() ImVec2

// Content boundaries max (e.g. window boundaries including scrolling, or current column boundaries). You should never need this. Always use GetCursorScreenPos() and GetContentRegionAvail()!
@[c:'ImGui_GetWindowContentRegionMin']
fn get_window_content_region_min() ImVec2

// Content boundaries min for the window (roughly (0,0)-Scroll), in window-local coordinates. You should never need this. Always use GetCursorScreenPos() and GetContentRegionAvail()!
@[c:'ImGui_GetWindowContentRegionMax']
fn get_window_content_region_max() ImVec2

// Content boundaries max for the window (roughly (0,0)+Size-Scroll), in window-local coordinates. You should never need this. Always use GetCursorScreenPos() and GetContentRegionAvail()!
// OBSOLETED in 1.90.0 (from September 2023)
@[c:'ImGui_BeginChildFrame']
fn begin_child_frame(id ID, size ImVec2) bool

// Implied window_flags = 0
@[c:'ImGui_BeginChildFrameEx']
fn begin_child_frame_ex(id ID, size ImVec2, window_flags WindowFlags) bool

@[c:'ImGui_EndChildFrame']
fn end_child_frame()

//static inline bool BeginChild(const char* str_id, const ImVec2& size_arg, bool borders, WindowFlags window_flags){ return BeginChild(str_id, size_arg, borders ? ChildFlags_Borders : ChildFlags_None, window_flags); } // Unnecessary as true == ChildFlags_Borders
//static inline bool BeginChild ID id, const ImVec2& size_arg, bool borders, WindowFlags window_flags)        { return BeginChild(id, size_arg, borders ? ChildFlags_Borders : ChildFlags_None, window_flags);     } // Unnecessary as true == ChildFlags_Borders
@[c:'ImGui_ShowStackToolWindow']
fn show_stack_tool_window(p_open &bool)

@[c:'ImGui_ComboObsolete']
fn combo_obsolete(label &i8, current_item &int, old_callback fn (voidptr, int, &&i8) bool, user_data voidptr, items_count int) bool

// Implied popup_max_height_in_items = -1
@[c:'ImGui_ComboObsoleteEx']
fn combo_obsolete_ex(label &i8, current_item &int, old_callback fn (voidptr, int, &&i8) bool, user_data voidptr, items_count int, popup_max_height_in_items int) bool

@[c:'ImGui_ListBoxObsolete']
fn list_box_obsolete(label &i8, current_item &int, old_callback fn (voidptr, int, &&i8) bool, user_data voidptr, items_count int) bool

// Implied height_in_items = -1
@[c:'ImGui_ListBoxObsoleteEx']
fn list_box_obsolete_ex(label &i8, current_item &int, old_callback fn (voidptr, int, &&i8) bool, user_data voidptr, items_count int, height_in_items int) bool

// OBSOLETED in 1.89.7 (from June 2023)
@[c:'ImGui_SetItemAllowOverlap']
fn set_item_allow_overlap()

// Use SetNextItemAllowOverlap() before item.
// OBSOLETED in 1.89.4 (from March 2023)
@[c:'ImGui_PushAllowKeyboardFocus']
fn push_allow_keyboard_focus(tab_stop bool)

@[c:'ImGui_PopAllowKeyboardFocus']
fn pop_allow_keyboard_focus()

// Some of the older obsolete names along with their replacement (commented out so they are not reported in IDE)
//-- OBSOLETED in 1.89 (from August 2022)
//IMGUI_API bool      ImageButton(ImTextureID user_texture_id, const ImVec2& size, const ImVec2& uv0 = ImVec2(0, 0), const ImVec2& uv1 = ImVec2(1, 1), int frame_padding = -1, const C.ImVec4& bg_col = C.ImVec4(0, 0, 0, 0), const C.ImVec4& tint_col = C.ImVec4(1, 1, 1, 1)); // --> Use new ImageButton() signature (explicit item id, regular FramePadding). Refer to code in 1.91 if you want to grab a copy of this version.
//-- OBSOLETED in 1.88 (from May 2022)
//static inline void  CaptureKeyboardFromApp(bool want_capture_keyboard = true)                   { SetNextFrameWantCaptureKeyboard(want_capture_keyboard); } // Renamed as name was misleading + removed default value.
//static inline void  CaptureMouseFromApp(bool want_capture_mouse = true)                         { SetNextFrameWantCaptureMouse(want_capture_mouse); }       // Renamed as name was misleading + removed default value.
//-- OBSOLETED in 1.87 (from February 2022, more formally obsoleted April 2024)
//IMGUI_API Key  GetKeyIndex Key key);                                                  { IM_ASSERT(key >= Key_NamedKey_BEGIN && key < Key_NamedKey_END); const ImGuiKeyData* key_data = GetKeyData(key); return  Key)(key_data - g.IO.KeysData); } // Map Key_* values into legacy native key index. == io.KeyMap[key]. When using a 1.87+ backend using io.AddKeyEvent(), calling GetKeyIndex() with ANY Key_XXXX values will return the same value!
//static inline Key GetKeyIndex Key key)                                                { IM_ASSERT(key >= Key_NamedKey_BEGIN && key < Key_NamedKey_END); return key; }
//-- OBSOLETED in 1.86 (from November 2021)
//IMGUI_API void      CalcListClipping(int items_count, float items_height, int* out_items_display_start, int* out_items_display_end); // Code removed, see 1.90 for last version of the code. Calculate range of visible items for large list of evenly sized items. Prefer using ImGuiListClipper.
//-- OBSOLETED in 1.85 (from August 2021)
//static inline float GetWindowContentRegionWidth()                                               { return GetWindowContentRegionMax().x - GetWindowContentRegionMin().x; }
//-- OBSOLETED in 1.81 (from February 2021)
//static inline bool  ListBoxHeader(const char* label, const ImVec2& size = ImVec2(0, 0))         { return BeginListBox(label, size); }
//static inline bool  ListBoxHeader(const char* label, int items_count, int height_in_items = -1) { float height = GetTextLineHeightWithSpacing() * ((height_in_items < 0 ? ImMin(items_count, 7) : height_in_items) + 0.25f) + GetStyle().FramePadding.y * 2.0f; return BeginListBox(label, ImVec2(0.0f, height)); } // Helper to calculate size from items_count and height_in_items
//static inline void  ListBoxFooter()                                                             { EndListBox(); }
//-- OBSOLETED in 1.79 (from August 2020)
//static inline void  OpenPopupContextItem(const char* str_id = NULL, MouseButton mb = 1)    { OpenPopupOnItemClick(str_id, mb); } // Bool return value removed. Use IsWindowAppearing() in BeginPopup() instead. Renamed in 1.77, renamed back in 1.79. Sorry!
//-- OBSOLETED in 1.78 (from June 2020): Old drag/sliders functions that took a 'float power > 1.0f' argument instead of SliderFlags_Logarithmic. See github.com/ocornut/imgui/issues/3361 for details.
//IMGUI_API bool      DragScalar(const char* label, DataType data_type, void* p_data, float v_speed, const void* p_min, const void* p_max, const char* format, float power = 1.0f)                                                            // OBSOLETED in 1.78 (from June 2020)
//IMGUI_API bool      DragScalarN(const char* label, DataType data_type, void* p_data, int components, float v_speed, const void* p_min, const void* p_max, const char* format, float power = 1.0f);                                          // OBSOLETED in 1.78 (from June 2020)
//IMGUI_API bool      SliderScalar(const char* label, DataType data_type, void* p_data, const void* p_min, const void* p_max, const char* format, float power = 1.0f);                                                                        // OBSOLETED in 1.78 (from June 2020)
//IMGUI_API bool      SliderScalarN(const char* label, DataType data_type, void* p_data, int components, const void* p_min, const void* p_max, const char* format, float power = 1.0f);                                                       // OBSOLETED in 1.78 (from June 2020)
//static inline bool  DragFloat(const char* label, float* v, float v_speed, float v_min, float v_max, const char* format, float power = 1.0f)    { return DragScalar(label, DataType_Float, v, v_speed, &v_min, &v_max, format, power); }     // OBSOLETED in 1.78 (from June 2020)
//static inline bool  DragFloat2(const char* label, float v[2], float v_speed, float v_min, float v_max, const char* format, float power = 1.0f) { return DragScalarN(label, DataType_Float, v, 2, v_speed, &v_min, &v_max, format, power); } // OBSOLETED in 1.78 (from June 2020)
//static inline bool  DragFloat3(const char* label, float v[3], float v_speed, float v_min, float v_max, const char* format, float power = 1.0f) { return DragScalarN(label, DataType_Float, v, 3, v_speed, &v_min, &v_max, format, power); } // OBSOLETED in 1.78 (from June 2020)
//static inline bool  DragFloat4(const char* label, float v[4], float v_speed, float v_min, float v_max, const char* format, float power = 1.0f) { return DragScalarN(label, DataType_Float, v, 4, v_speed, &v_min, &v_max, format, power); } // OBSOLETED in 1.78 (from June 2020)
//static inline bool  SliderFloat(const char* label, float* v, float v_min, float v_max, const char* format, float power = 1.0f)                 { return SliderScalar(label, DataType_Float, v, &v_min, &v_max, format, power); }            // OBSOLETED in 1.78 (from June 2020)
//static inline bool  SliderFloat2(const char* label, float v[2], float v_min, float v_max, const char* format, float power = 1.0f)              { return SliderScalarN(label, DataType_Float, v, 2, &v_min, &v_max, format, power); }        // OBSOLETED in 1.78 (from June 2020)
//static inline bool  SliderFloat3(const char* label, float v[3], float v_min, float v_max, const char* format, float power = 1.0f)              { return SliderScalarN(label, DataType_Float, v, 3, &v_min, &v_max, format, power); }        // OBSOLETED in 1.78 (from June 2020)
//static inline bool  SliderFloat4(const char* label, float v[4], float v_min, float v_max, const char* format, float power = 1.0f)              { return SliderScalarN(label, DataType_Float, v, 4, &v_min, &v_max, format, power); }        // OBSOLETED in 1.78 (from June 2020)
//-- OBSOLETED in 1.77 and before
//static inline bool  BeginPopupContextWindow(const char* str_id, MouseButton mb, bool over_items) { return BeginPopupContextWindow(str_id, mb | (over_items ? 0 : PopupFlags_NoOpenOverItems)); } // OBSOLETED in 1.77 (from June 2020)
//static inline void  TreeAdvanceToLabelPos()               { SetCursorPosX(GetCursorPosX() + GetTreeNodeToLabelSpacing()); }   // OBSOLETED in 1.72 (from July 2019)
//static inline void  SetNextTreeNodeOpen(bool open, Cond cond = 0) { SetNextItemOpen(open, cond); }                       // OBSOLETED in 1.71 (from June 2019)
//static inline float GetContentRegionAvailWidth()          { return GetContentRegionAvail().x; }                               // OBSOLETED in 1.70 (from May 2019)
//static inline ImDrawList* GetOverlayDrawList()            { return GetForegroundDrawList(); }                                 // OBSOLETED in 1.69 (from Mar 2019)
//static inline void  SetScrollHere(float ratio = 0.5f)     { SetScrollHereY(ratio); }                                          // OBSOLETED in 1.66 (from Nov 2018)
//static inline bool  IsItemDeactivatedAfterChange()        { return IsItemDeactivatedAfterEdit(); }                            // OBSOLETED in 1.63 (from Aug 2018)
//-- OBSOLETED in 1.60 and before
//static inline bool  IsAnyWindowFocused()                  { return IsWindowFocused FocusedFlags_AnyWindow); }            // OBSOLETED in 1.60 (from Apr 2018)
//static inline bool  IsAnyWindowHovered()                  { return IsWindowHovered HoveredFlags_AnyWindow); }            // OBSOLETED in 1.60 (between Dec 2017 and Apr 2018)
//static inline void  ShowTestWindow()                      { return ShowDemoWindow(); }                                        // OBSOLETED in 1.53 (between Oct 2017 and Dec 2017)
//static inline bool  IsRootWindowFocused()                 { return IsWindowFocused FocusedFlags_RootWindow); }           // OBSOLETED in 1.53 (between Oct 2017 and Dec 2017)
//static inline bool  IsRootWindowOrAnyChildFocused()       { return IsWindowFocused FocusedFlags_RootAndChildWindows); }  // OBSOLETED in 1.53 (between Oct 2017 and Dec 2017)
//static inline void  SetNextWindowContentWidth(float w)    { SetNextWindowContentSize(ImVec2(w, 0.0f)); }                      // OBSOLETED in 1.53 (between Oct 2017 and Dec 2017)
//static inline float GetItemsLineHeightWithSpacing()       { return GetFrameHeightWithSpacing(); }                             // OBSOLETED in 1.53 (between Oct 2017 and Dec 2017)
//IMGUI_API bool      Begin(char* name, bool* p_open, ImVec2 size_first_use, float bg_alpha = -1.0f, WindowFlags flags=0); // OBSOLETED in 1.52 (between Aug 2017 and Oct 2017): Equivalent of using SetNextWindowSize(size, Cond_FirstUseEver) and SetNextWindowBgAlpha().
//static inline bool  IsRootWindowOrAnyChildHovered()       { return IsWindowHovered HoveredFlags_RootAndChildWindows); }  // OBSOLETED in 1.52 (between Aug 2017 and Oct 2017)
//static inline void  AlignFirstTextHeightToWidgets()       { AlignTextToFramePadding(); }                                      // OBSOLETED in 1.52 (between Aug 2017 and Oct 2017)
//static inline void  SetNextWindowPosCenter Cond c=0) { SetNextWindowPos(GetMainViewport()->GetCenter(), c, ImVec2(0.5f,0.5f)); } // OBSOLETED in 1.52 (between Aug 2017 and Oct 2017)
//static inline bool  IsItemHoveredRect()                   { return IsItemHovered HoveredFlags_RectOnly); }               // OBSOLETED in 1.51 (between Jun 2017 and Aug 2017)
//static inline bool  IsPosHoveringAnyWindow(const ImVec2&) { IM_ASSERT(0); return false; }                                     // OBSOLETED in 1.51 (between Jun 2017 and Aug 2017): This was misleading and partly broken. You probably want to use the io.WantCaptureMouse flag instead.
//static inline bool  IsMouseHoveringAnyWindow()            { return IsWindowHovered HoveredFlags_AnyWindow); }            // OBSOLETED in 1.51 (between Jun 2017 and Aug 2017)
//static inline bool  IsMouseHoveringWindow()               { return IsWindowHovered HoveredFlags_AllowWhenBlockedByPopup | HoveredFlags_AllowWhenBlockedByActiveItem); }       // OBSOLETED in 1.51 (between Jun 2017 and Aug 2017)
//-- OBSOLETED in 1.50 and before
//static inline bool  CollapsingHeader(char* label, const char* str_id, bool framed = true, bool default_open = false) { return CollapsingHeader(label, (default_open ? (1 << 5) : 0)); } // OBSOLETED in 1.49
//static inline ImFont*GetWindowFont()                      { return GetFont(); }                                               // OBSOLETED in 1.48
//static inline float GetWindowFontSize()                   { return GetFontSize(); }                                           // OBSOLETED in 1.48
//static inline void  SetScrollPosHere()                    { SetScrollHere(); }                                                // OBSOLETED in 1.42
//-- OBSOLETED in 1.82 (from Mars 2021): flags for AddRect(), AddRectFilled(), AddImageRounded(), PathRect()
//typedef ImDrawFlags ImDrawCornerFlags;
//enum ImDrawCornerFlags_
//{
//    ImDrawCornerFlags_None      = ImDrawFlags_RoundCornersNone,         // Was == 0 prior to 1.82, this is now == ImDrawFlags_RoundCornersNone which is != 0 and not implicit
//    ImDrawCornerFlags_TopLeft   = ImDrawFlags_RoundCornersTopLeft,      // Was == 0x01 (1 << 0) prior to 1.82. Order matches ImDrawFlags_NoRoundCorner* flag (we exploit this internally).
//    ImDrawCornerFlags_TopRight  = ImDrawFlags_RoundCornersTopRight,     // Was == 0x02 (1 << 1) prior to 1.82.
//    ImDrawCornerFlags_BotLeft   = ImDrawFlags_RoundCornersBottomLeft,   // Was == 0x04 (1 << 2) prior to 1.82.
//    ImDrawCornerFlags_BotRight  = ImDrawFlags_RoundCornersBottomRight,  // Was == 0x08 (1 << 3) prior to 1.82.
//    ImDrawCornerFlags_All       = ImDrawFlags_RoundCornersAll,          // Was == 0x0F prior to 1.82
//    ImDrawCornerFlags_Top       = ImDrawCornerFlags_TopLeft | ImDrawCornerFlags_TopRight,
//    ImDrawCornerFlags_Bot       = ImDrawCornerFlags_BotLeft | ImDrawCornerFlags_BotRight,
//    ImDrawCornerFlags_Left      = ImDrawCornerFlags_TopLeft | ImDrawCornerFlags_BotLeft,
//    ImDrawCornerFlags_Right     = ImDrawCornerFlags_TopRight | ImDrawCornerFlags_BotRight,
//};
// RENAMED and MERGED both Key_ModXXX and ModFlags_XXX into Mod_XXX (from September 2022)
// RENAMED KeyModFlags -> ModFlags in 1.88 (from April 2022). Exceptionally commented out ahead of obscolescence schedule to reduce confusion and because they were not meant to be used in the first place.
//typedef KeyChord ModFlags;      // == int. We generally use KeyChord to mean "a Key or-ed with any number of Mod_XXX value", so you may store mods in there.
//enum ModFlags_ { ModFlags_None = 0, ModFlags_Ctrl = Mod_Ctrl, ModFlags_Shift = Mod_Shift, ModFlags_Alt = Mod_Alt, ModFlags_Super = Mod_Super };
//typedef KeyChord KeyModFlags; // == int
//enum KeyModFlags_ { KeyModFlags_None = 0, KeyModFlags_Ctrl = Mod_Ctrl, KeyModFlags_Shift = Mod_Shift, KeyModFlags_Alt = Mod_Alt, KeyModFlags_Super = Mod_Super };
// OBSOLETED IN 1.90 (now using C++11 standard version)
// #ifndef IMGUI_DISABLE_OBSOLETE_FUNCTIONS
// RENAMED IMGUI_DISABLE_METRICS_WINDOW > IMGUI_DISABLE_DEBUG_TOOLS in 1.88 (from June 2022)
// #ifdef IMGUI_DISABLE_METRICS_WINDOW
//-----------------------------------------------------------------------------
// #if defined(__GNUC__)
// #if defined(__clang__)
// #ifdef _MSC_VER
// Include imgui_user.h at the end of imgui.h
// May be convenient for some users to only explicitly include vanilla imgui.h and have extra stuff included.
// #ifdef IMGUI_USER_H_FILENAME
// #ifdef IMGUI_INCLUDE_IMGUI_USER_H
// #ifndef IMGUI_DISABLE
// End of extern "C" block
