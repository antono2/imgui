module imgui


#flag -I @VMODROOT/include
#flag -I @VMODROOT/include/imgui
#flag -I @VMODROOT/include/imgui/backends
#flag @VMODROOT/lib/libcimgui.so

#define CIMGUI_DEFINE_ENUMS_AND_STRUCTS
#define IMGUI_USE_WCHAR32

#include "cimgui.h"

