@[translated]
module imgui


pub const version = "1.91.9b"
pub const version_num = 19191

pub type DockNodeSettings = C.ImGuiDockNodeSettings
@[typedef]
pub struct C.ImGuiDockNodeSettings {}

pub type SizeCallback = fn(&SizeCallbackData)
pub type TextFilter = C.ImGuiTextFilter
@[typedef]
pub struct C.ImGuiTextFilter {
pub mut:
  InputBuf [256]char
  Filters ImVector_TextRange
  CountGrep int
}
pub type Va_list = C.va_list
@[typedef]
pub struct C.va_list {}

pub type InputTextCallback = fn(&InputTextCallbackData) int

pub type ImWchar = u32
pub type DockRequest = C.ImGuiDockRequest
@[typedef]
pub struct C.ImGuiDockRequest {}

// This file is automatically generated by generator.lua from https://github.com/cimgui/cimgui
// based on imgui.h file version "1.91.9b" 19191 from Dear ImGui https://github.com/ocornut/imgui
// with imgui_internal.h api
// with imgui_freetype.h api
// docking branch
// typedef unsigned long long ImU64;


pub type ImVector_const_charPtr = C.ImVector_const_charPtr
@[typedef]
struct C.ImVector_const_charPtr {
pub mut:
	Size     int
	Capacity int
	Data     /*&&u8*/voidptr= unsafe{ nil }
}

type ID = u32
type ImS8 = i8
type ImU8 = u8
type ImS16 = i16
type ImU16 = u16
type ImS32 = int
type ImU32 = u32
type ImS64 = i64
type ImU64 = i64
type Col = int
type Cond = int
type DataType = int
type MouseButton = int
type MouseCursor = int
type StyleVar = int
type TableBgTarget = int
type ImDrawFlags = int
type ImDrawListFlags = int
type ImFontAtlasFlags = int
type BackendFlags = int
type ButtonFlags = int
type ChildFlags = int
type ColorEditFlags = int
type ConfigFlags = int
type ComboFlags = int
type DockNodeFlags = int
type DragDropFlags = int
type FocusedFlags = int
type HoveredFlags = int
type InputFlags = int
type InputTextFlags = int
type ItemFlags = int
type KeyChord = int
type PopupFlags = int
type MultiSelectFlags = int
type SelectableFlags = int
type SliderFlags = int
type TabBarFlags = int
type TabItemFlags = int
type TableFlags = int
type TableColumnFlags = int
type TableRowFlags = int
type TreeNodeFlags = int
type ViewportFlags = int
type WindowFlags = int
type ImWchar32 = u32
type ImWchar16 = u16
type SelectionUserData = i64
type MemAllocFunc = fn (usize, voidptr) voidptr

type MemFreeFunc = fn (voidptr, voidptr)



pub type ImVec2 = C.ImVec2
@[typedef]
struct C.ImVec2 {
pub mut:

	x f32
	y f32
}



pub type ImVec4 = C.ImVec4
@[typedef]
struct C.ImVec4 {
pub mut:

	x f32
	y f32
	z f32
	w f32
}

type ImTextureID = i64

enum WindowFlags_ {
 none                        = 0
 no_title_bar                = 1 << 0
 no_resize                   = 1 << 1
 no_move                     = 1 << 2
 no_scrollbar                = 1 << 3
 no_scroll_with_mouse        = 1 << 4
 no_collapse                 = 1 << 5
 always_auto_resize          = 1 << 6
 no_background               = 1 << 7
 no_saved_settings           = 1 << 8
 no_mouse_inputs             = 1 << 9
 menu_bar                    = 1 << 10
 horizontal_scrollbar        = 1 << 11
 no_focus_on_appearing       = 1 << 12
 no_bring_to_front_on_focus  = 1 << 13
 always_vertical_scrollbar   = 1 << 14
 always_horizontal_scrollbar = 1 << 15
 no_nav_inputs               = 1 << 16
 no_nav_focus                = 1 << 17
 unsaved_document            = 1 << 18
 no_docking                  = 1 << 19
 no_nav                      = 1 << 16 | 1 << 17
 no_decoration               = 1 << 0 | 1 << 1 | 1 << 3 | 1 << 5
 no_inputs                   = 1 << 9 | 1 << 16 | 1 << 17
 dock_node_host              = 1 << 23
 child_window                = 1 << 24
 tooltip                     = 1 << 25
 popup                       = 1 << 26
 modal                       = 1 << 27
 child_menu                  = 1 << 28
}

enum ChildFlags_ {
 none                      = 0
 borders                   = 1 << 0
 always_use_window_padding = 1 << 1
 resize_x                  = 1 << 2
 resize_y                  = 1 << 3
 auto_resize_x             = 1 << 4
 auto_resize_y             = 1 << 5
 always_auto_resize        = 1 << 6
 frame_style               = 1 << 7
 nav_flattened             = 1 << 8
}

enum ItemFlags_ {
 none                 = 0
 no_tab_stop          = 1 << 0
 no_nav               = 1 << 1
 no_nav_default_focus = 1 << 2
 button_repeat        = 1 << 3
 auto_close_popups    = 1 << 4
 allow_duplicate_id   = 1 << 5
}

enum InputTextFlags_ {
 none                    = 0
 chars_decimal           = 1 << 0
 chars_hexadecimal       = 1 << 1
 chars_scientific        = 1 << 2
 chars_uppercase         = 1 << 3
 chars_no_blank          = 1 << 4
 allow_tab_input         = 1 << 5
 enter_returns_true      = 1 << 6
 escape_clears_all       = 1 << 7
 ctrl_enter_for_new_line = 1 << 8
 read_only               = 1 << 9
 password                = 1 << 10
 always_overwrite        = 1 << 11
 auto_select_all         = 1 << 12
 parse_empty_ref_val     = 1 << 13
 display_empty_ref_val   = 1 << 14
 no_horizontal_scroll    = 1 << 15
 no_undo_redo            = 1 << 16
 elide_left              = 1 << 17
 callback_completion     = 1 << 18
 callback_history        = 1 << 19
 callback_always         = 1 << 20
 callback_char_filter    = 1 << 21
 callback_resize         = 1 << 22
 callback_edit           = 1 << 23
}

enum TreeNodeFlags_ {
 none                     = 0
 selected                 = 1 << 0
 framed                   = 1 << 1
 allow_overlap            = 1 << 2
 no_tree_push_on_open     = 1 << 3
 no_auto_open_on_log      = 1 << 4
 default_open             = 1 << 5
 open_on_double_click     = 1 << 6
 open_on_arrow            = 1 << 7
 leaf                     = 1 << 8
 bullet                   = 1 << 9
 frame_padding            = 1 << 10
 span_avail_width         = 1 << 11
 span_full_width          = 1 << 12
 span_label_width         = 1 << 13
 span_all_columns         = 1 << 14
 label_span_all_columns   = 1 << 15
 nav_left_jumps_back_here = 1 << 17
 collapsing_header        = 1 << 1 | 1 << 3 | 1 << 4
}

enum PopupFlags_ {
 //none                        = 0
 mouse_button_left           = 0
 mouse_button_right          = 1
 mouse_button_middle         = 2
 mouse_button_mask_          = 31
 //mouse_button_default_       = 1
 no_reopen                   = 1 << 5
 no_open_over_existing_popup = 1 << 7
 no_open_over_items          = 1 << 8
 any_popup_id                = 1 << 10
 any_popup_level             = 1 << 11
 any_popup                   = 1 << 10 | 1 << 11
}

enum SelectableFlags_ {
 none                 = 0
 no_auto_close_popups = 1 << 0
 span_all_columns     = 1 << 1
 allow_double_click   = 1 << 2
 disabled             = 1 << 3
 allow_overlap        = 1 << 4
 highlight            = 1 << 5
}

enum ComboFlags_ {
 none              = 0
 popup_align_left  = 1 << 0
 height_small      = 1 << 1
 height_regular    = 1 << 2
 height_large      = 1 << 3
 height_largest    = 1 << 4
 no_arrow_button   = 1 << 5
 no_preview        = 1 << 6
 width_fit_preview = 1 << 7
 height_mask_      = 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4
}

enum TabBarFlags_ {
 none                              = 0
 reorderable                       = 1 << 0
 auto_select_new_tabs              = 1 << 1
 tab_list_popup_button             = 1 << 2
 no_close_with_middle_mouse_button = 1 << 3
 no_tab_list_scrolling_buttons     = 1 << 4
 no_tooltip                        = 1 << 5
 draw_selected_overline            = 1 << 6
 fitting_policy_resize_down        = 1 << 7
 fitting_policy_scroll             = 1 << 8
 fitting_policy_mask_              = 1 << 7 | 1 << 8
 //fitting_policy_default_           = 1 << 7
}

enum TabItemFlags_ {
 none                              = 0
 unsaved_document                  = 1 << 0
 set_selected                      = 1 << 1
 no_close_with_middle_mouse_button = 1 << 2
 no_push_id                        = 1 << 3
 no_tooltip                        = 1 << 4
 no_reorder                        = 1 << 5
 leading                           = 1 << 6
 trailing                          = 1 << 7
 no_assumed_closure                = 1 << 8
}

enum FocusedFlags_ {
 none                   = 0
 child_windows          = 1 << 0
 root_window            = 1 << 1
 any_window             = 1 << 2
 no_popup_hierarchy     = 1 << 3
 dock_hierarchy         = 1 << 4
 root_and_child_windows = 1 << 1 | 1 << 0
}

enum HoveredFlags_ {
 none                              = 0
 child_windows                     = 1 << 0
 root_window                       = 1 << 1
 any_window                        = 1 << 2
 no_popup_hierarchy                = 1 << 3
 dock_hierarchy                    = 1 << 4
 allow_when_blocked_by_popup       = 1 << 5
 allow_when_blocked_by_active_item = 1 << 7
 allow_when_overlapped_by_item     = 1 << 8
 allow_when_overlapped_by_window   = 1 << 9
 allow_when_disabled               = 1 << 10
 no_nav_override                   = 1 << 11
 allow_when_overlapped             = 1 << 8 | 1 << 9
 rect_only                         = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9
 root_and_child_windows            = 1 << 1 | 1 << 0
 for_tooltip                       = 1 << 12
 stationary                        = 1 << 13
 delay_none                        = 1 << 14
 delay_short                       = 1 << 15
 delay_normal                      = 1 << 16
 no_shared_delay                   = 1 << 17
}

enum DockNodeFlags_ {
 none                         = 0
 keep_alive_only              = 1 << 0
 no_docking_over_central_node = 1 << 2
 passthru_central_node        = 1 << 3
 no_docking_split             = 1 << 4
 no_resize                    = 1 << 5
 auto_hide_tab_bar            = 1 << 6
 no_undocking                 = 1 << 7
}

enum DragDropFlags_ {
 none                          = 0
 source_no_preview_tooltip     = 1 << 0
 source_no_disable_hover       = 1 << 1
 source_no_hold_to_open_others = 1 << 2
 source_allow_null_id          = 1 << 3
 source_extern                 = 1 << 4
 payload_auto_expire           = 1 << 5
 payload_no_cross_context      = 1 << 6
 payload_no_cross_process      = 1 << 7
 accept_before_delivery        = 1 << 10
 accept_no_draw_default_rect   = 1 << 11
 accept_no_preview_tooltip     = 1 << 12
 accept_peek_only              = 1 << 10 | 1 << 11
}

enum DataType_ {
 s8
 u8
 s16
 u16
 s32
 u32
 s64
 u64
 float
 double
 bool
 string
 count
}

enum Dir {
 none  = -1
 left  = 0
 right = 1
 up    = 2
 down  = 3
 count = 4
}

enum SortDirection {
 none       = 0
 ascending  = 1
 descending = 2
}

enum Key {
 none                   = 0
//named_begin        = 512
 tab                    = 512
 left_arrow             = 513
 right_arrow            = 514
 up_arrow               = 515
 down_arrow             = 516
 page_up                = 517
 page_down              = 518
 home                   = 519
 end                    = 520
 insert                 = 521
 delete                 = 522
 backspace              = 523
 space                  = 524
 enter                  = 525
 escape                 = 526
 left_ctrl              = 527
 left_shift             = 528
 left_alt               = 529
 left_super             = 530
 right_ctrl             = 531
 right_shift            = 532
 right_alt              = 533
 right_super            = 534
 menu                   = 535
 _0 = 536
 _1 = 537
 _2 = 538
 _3 = 539
 _4 = 540
 _5 = 541
 _6 = 542
 _7 = 543
 _8 = 544
 _9 = 545
 a                      = 546
 b                      = 547
 c                      = 548
 d                      = 549
 e                      = 550
 f                      = 551
 g                      = 552
 h                      = 553
 i                      = 554
 j                      = 555
 k                      = 556
 l                      = 557
 m                      = 558
 n                      = 559
 o                      = 560
 p                      = 561
 q                      = 562
 r                      = 563
 s                      = 564
 t                      = 565
 u                      = 566
 v                      = 567
 w                      = 568
 x                      = 569
 y                      = 570
 z                      = 571
 f1                     = 572
 f2                     = 573
 f3                     = 574
 f4                     = 575
 f5                     = 576
 f6                     = 577
 f7                     = 578
 f8                     = 579
 f9                     = 580
 f10                    = 581
 f11                    = 582
 f12                    = 583
 f13                    = 584
 f14                    = 585
 f15                    = 586
 f16                    = 587
 f17                    = 588
 f18                    = 589
 f19                    = 590
 f20                    = 591
 f21                    = 592
 f22                    = 593
 f23                    = 594
 f24                    = 595
 apostrophe             = 596
 comma                  = 597
 minus                  = 598
 period                 = 599
 slash                  = 600
 semicolon              = 601
 equal                  = 602
 left_bracket           = 603
 backslash              = 604
 right_bracket          = 605
 grave_accent           = 606
 caps_lock              = 607
 scroll_lock            = 608
 num_lock               = 609
 print_screen           = 610
 pause                  = 611
 pad0                = 612
 pad1                = 613
 pad2                = 614
 pad3                = 615
 pad4                = 616
 pad5                = 617
 pad6                = 618
 pad7                = 619
 pad8                = 620
 pad9                = 621
 pad_decimal         = 622
 pad_divide          = 623
 pad_multiply        = 624
 pad_subtract        = 625
 pad_add             = 626
 pad_enter           = 627
 pad_equal           = 628
 app_back               = 629
 app_forward            = 630
 oem102                 = 631
 gamepad_start          = 632
 gamepad_back           = 633
 gamepad_face_left      = 634
 gamepad_face_right     = 635
 gamepad_face_up        = 636
 gamepad_face_down      = 637
 gamepad_dpad_left      = 638
 gamepad_dpad_right     = 639
 gamepad_dpad_up        = 640
 gamepad_dpad_down      = 641
 gamepad_l1             = 642
 gamepad_r1             = 643
 gamepad_l2             = 644
 gamepad_r2             = 645
 gamepad_l3             = 646
 gamepad_r3             = 647
 gamepad_ls_tick_left   = 648
 gamepad_ls_tick_right  = 649
 gamepad_ls_tick_up     = 650
 gamepad_ls_tick_down   = 651
 gamepad_rs_tick_left   = 652
 gamepad_rs_tick_right  = 653
 gamepad_rs_tick_up     = 654
 gamepad_rs_tick_down   = 655
 mouse_left             = 656
 mouse_right            = 657
 mouse_middle           = 658
 mouse_x1               = 659
 mouse_x2               = 660
 mouse_wheel_x          = 661
 mouse_wheel_y          = 662
 reserved_for_mod_ctrl  = 663
 reserved_for_mod_shift = 664
 reserved_for_mod_alt   = 665
 reserved_for_mod_super = 666
 named_end          = 667
//mod_none                   = 0
 mod_ctrl                   = 1 << 12
 mod_shift                  = 1 << 13
 mod_alt                    = 1 << 14
 mod_super                  = 1 << 15
 mod_mask_                  = 61440
 named_count        = 667 - 512
}

enum InputFlags_ {
 none                    = 0
 repeat                  = 1 << 0
 route_active            = 1 << 10
 route_focused           = 1 << 11
 route_global            = 1 << 12
 route_always            = 1 << 13
 route_over_focused      = 1 << 14
 route_over_active       = 1 << 15
 route_unless_bg_focused = 1 << 16
 route_from_root_window  = 1 << 17
 tooltip                 = 1 << 18
}

enum ConfigFlags_ {
 none                       = 0
 nav_enable_keyboard        = 1 << 0
 nav_enable_gamepad         = 1 << 1
 no_mouse                   = 1 << 4
 no_mouse_cursor_change     = 1 << 5
 no_keyboard                = 1 << 6
 docking_enable             = 1 << 7
 viewports_enable           = 1 << 10
 dpi_enable_scale_viewports = 1 << 14
 dpi_enable_scale_fonts     = 1 << 15
 is_srgb                    = 1 << 20
 is_touch_screen            = 1 << 21
}

enum BackendFlags_ {
 none                       = 0
 has_gamepad                = 1 << 0
 has_mouse_cursors          = 1 << 1
 has_set_mouse_pos          = 1 << 2
 renderer_has_vtx_offset    = 1 << 3
 platform_has_viewports     = 1 << 10
 has_mouse_hovered_viewport = 1 << 11
 renderer_has_viewports     = 1 << 12
}

enum Col_ {
 text
 text_disabled
 window_bg
 child_bg
 popup_bg
 border
 border_shadow
 frame_bg
 frame_bg_hovered
 frame_bg_active
 title_bg
 title_bg_active
 title_bg_collapsed
 menu_bar_bg
 scrollbar_bg
 scrollbar_grab
 scrollbar_grab_hovered
 scrollbar_grab_active
 check_mark
 slider_grab
 slider_grab_active
 button
 button_hovered
 button_active
 header
 header_hovered
 header_active
 separator
 separator_hovered
 separator_active
 resize_grip
 resize_grip_hovered
 resize_grip_active
 tab_hovered
 tab
 tab_selected
 tab_selected_overline
 tab_dimmed
 tab_dimmed_selected
 tab_dimmed_selected_overline
 docking_preview
 docking_empty_bg
 plot_lines
 plot_lines_hovered
 plot_histogram
 plot_histogram_hovered
 table_header_bg
 table_border_strong
 table_border_light
 table_row_bg
 table_row_bg_alt
 text_link
 text_selected_bg
 drag_drop_target
 nav_cursor
 nav_windowing_highlight
 nav_windowing_dim_bg
 modal_window_dim_bg
 count
}

enum StyleVar_ {
 alpha
 disabled_alpha
 window_padding
 window_rounding
 window_border_size
 window_min_size
 window_title_align
 child_rounding
 child_border_size
 popup_rounding
 popup_border_size
 frame_padding
 frame_rounding
 frame_border_size
 item_spacing
 item_inner_spacing
 indent_spacing
 cell_padding
 scrollbar_size
 scrollbar_rounding
 grab_min_size
 grab_rounding
 image_border_size
 tab_rounding
 tab_border_size
 tab_bar_border_size
 tab_bar_overline_size
 table_angled_headers_angle
 table_angled_headers_text_align
 button_text_align
 selectable_text_align
 separator_text_border_size
 separator_text_align
 separator_text_padding
 docking_separator_size
 count
}

enum ButtonFlags_ {
 none                = 0
 mouse_button_left   = 1 << 0
 mouse_button_right  = 1 << 1
 mouse_button_middle = 1 << 2
 mouse_button_mask_  = 1 << 0 | 1 << 1 | 1 << 2
 enable_nav          = 1 << 3
}

enum ColorEditFlags_ {
 none               = 0
 no_alpha           = 1 << 1
 no_picker          = 1 << 2
 no_options         = 1 << 3
 no_small_preview   = 1 << 4
 no_inputs          = 1 << 5
 no_tooltip         = 1 << 6
 no_label           = 1 << 7
 no_side_preview    = 1 << 8
 no_drag_drop       = 1 << 9
 no_border          = 1 << 10
 alpha_opaque       = 1 << 11
 alpha_no_bg        = 1 << 12
 alpha_preview_half = 1 << 13
 alpha_bar          = 1 << 16
 hdr                = 1 << 19
 display_rgb        = 1 << 20
 display_hsv        = 1 << 21
 display_hex        = 1 << 22
 uint8              = 1 << 23
 float              = 1 << 24
 picker_hue_bar     = 1 << 25
 picker_hue_wheel   = 1 << 26
 input_rgb          = 1 << 27
 input_hsv          = 1 << 28
 default_options_   = 1 << 23 | 1 << 20 | 1 << 27 | 1 << 25
 alpha_mask_        = 1 << 1 | 1 << 11 | 1 << 12 | 1 << 13
 display_mask_      = 1 << 20 | 1 << 21 | 1 << 22
 data_type_mask_    = 1 << 23 | 1 << 24
 picker_mask_       = 1 << 26 | 1 << 25
 input_mask_        = 1 << 27 | 1 << 28
}

enum SliderFlags_ {
 none               = 0
 logarithmic        = 1 << 5
 no_round_to_format = 1 << 6
 no_input           = 1 << 7
 wrap_around        = 1 << 8
 clamp_on_input     = 1 << 9
 clamp_zero_range   = 1 << 10
 no_speed_tweaks    = 1 << 11
 always_clamp       = 1 << 9 | 1 << 10
 invalid_mask_      = 1879048207
}

enum MouseButton_ {
 left   = 0
 right  = 1
 middle = 2
 count  = 5
}

enum MouseCursor_ {
 none  = -1
 arrow = 0
 text_input
 resize_all
 resize_ns
 resize_ew
 resize_nesw
 resize_nwse
 hand
 wait
 progress
 not_allowed
 count
}

enum MouseSource {
 mouse        = 0
 touch_screen = 1
 pen          = 2
 count        = 3
}

enum Cond_ {
 none           = 0
 always         = 1 << 0
 once           = 1 << 1
 first_use_ever = 1 << 2
 appearing      = 1 << 3
}

enum TableFlags_ {
 none                            = 0
 resizable                       = 1 << 0
 reorderable                     = 1 << 1
 hideable                        = 1 << 2
 sortable                        = 1 << 3
 no_saved_settings               = 1 << 4
 context_menu_in_body            = 1 << 5
 row_bg                          = 1 << 6
 borders_inner_h                 = 1 << 7
 borders_outer_h                 = 1 << 8
 borders_inner_v                 = 1 << 9
 borders_outer_v                 = 1 << 10
 borders_h                       = 1 << 7 | 1 << 8
 borders_v                       = 1 << 9 | 1 << 10
 borders_inner                   = 1 << 9 | 1 << 7
 borders_outer                   = 1 << 10 | 1 << 8
 borders                         = 1 << 9 | 1 << 7 | 1 << 10 | 1 << 8
 no_borders_in_body              = 1 << 11
 no_borders_in_body_until_resize = 1 << 12
 sizing_fixed_fit                = 1 << 13
 sizing_fixed_same               = 2 << 13
 sizing_stretch_prop             = 3 << 13
 sizing_stretch_same             = 4 << 13
 no_host_extend_x                = 1 << 16
 no_host_extend_y                = 1 << 17
 no_keep_columns_visible         = 1 << 18
 precise_widths                  = 1 << 19
 no_clip                         = 1 << 20
 pad_outer_x                     = 1 << 21
 no_pad_outer_x                  = 1 << 22
 no_pad_inner_x                  = 1 << 23
 scroll_x                        = 1 << 24
 scroll_y                        = 1 << 25
 sort_multi                      = 1 << 26
 sort_tristate                   = 1 << 27
 highlight_hovered_column        = 1 << 28
 sizing_mask_                    = 1 << 13 | 2 << 13 | 3 << 13 | 4 << 13
}

enum TableColumnFlags_ {
 none                   = 0
 disabled               = 1 << 0
 default_hide           = 1 << 1
 default_sort           = 1 << 2
 width_stretch          = 1 << 3
 width_fixed            = 1 << 4
 no_resize              = 1 << 5
 no_reorder             = 1 << 6
 no_hide                = 1 << 7
 no_clip                = 1 << 8
 no_sort                = 1 << 9
 no_sort_ascending      = 1 << 10
 no_sort_descending     = 1 << 11
 no_header_label        = 1 << 12
 no_header_width        = 1 << 13
 prefer_sort_ascending  = 1 << 14
 prefer_sort_descending = 1 << 15
 indent_enable          = 1 << 16
 indent_disable         = 1 << 17
 angled_header          = 1 << 18
 is_enabled             = 1 << 24
 is_visible             = 1 << 25
 is_sorted              = 1 << 26
 is_hovered             = 1 << 27
 width_mask_            = 1 << 3 | 1 << 4
 indent_mask_           = 1 << 16 | 1 << 17
 status_mask_           = 1 << 24 | 1 << 25 | 1 << 26 | 1 << 27
 no_direct_resize_      = 1 << 30
}

enum TableRowFlags_ {
 none    = 0
 headers = 1 << 0
}

enum TableBgTarget_ {
 none    = 0
 row_bg0 = 1
 row_bg1 = 2
 cell_bg = 3
}



pub type TableSortSpecs = C.ImGuiTableSortSpecs
@[typedef]
struct C.ImGuiTableSortSpecs {
pub mut:
	Specs      /*&TableColumnSortSpecs*/voidptr= unsafe{ nil }
	SpecsCount int
	SpecsDirty bool
}



pub type TableColumnSortSpecs = C.ImGuiTableColumnSortSpecs
@[typedef]
struct C.ImGuiTableColumnSortSpecs {
pub mut:
	ColumnUserID  ID
	ColumnIndex   ImS16
	SortOrder     ImS16
	SortDirection SortDirection
}



pub type Style = C.ImGuiStyle
@[typedef]
struct C.ImGuiStyle {
pub mut:
	Alpha                            f32
	DisabledAlpha                    f32
	WindowPadding                    ImVec2
	WindowRounding                   f32
	WindowBorderSize                 f32
	WindowBorderHoverPadding         f32
	WindowMinSize                    ImVec2
	WindowTitleAlign                 ImVec2
	WindowMenuButtonPosition         Dir
	ChildRounding                    f32
	ChildBorderSize                  f32
	PopupRounding                    f32
	PopupBorderSize                  f32
	FramePadding                     ImVec2
	FrameRounding                    f32
	FrameBorderSize                  f32
	ItemSpacing                      ImVec2
	ItemInnerSpacing                 ImVec2
	CellPadding                      ImVec2
	TouchExtraPadding                ImVec2
	IndentSpacing                    f32
	ColumnsMinSpacing                f32
	ScrollbarSize                    f32
	ScrollbarRounding                f32
	GrabMinSize                      f32
	GrabRounding                     f32
	LogSliderDeadzone                f32
	ImageBorderSize                  f32
	TabRounding                      f32
	TabBorderSize                    f32
	TabCloseButtonMinWidthSelected   f32
	TabCloseButtonMinWidthUnselected f32
	TabBarBorderSize                 f32
	TabBarOverlineSize               f32
	TableAngledHeadersAngle          f32
	TableAngledHeadersTextAlign      ImVec2
	ColorButtonPosition              Dir
	ButtonTextAlign                  ImVec2
	SelectableTextAlign              ImVec2
	SeparatorTextBorderSize          f32
	SeparatorTextAlign               ImVec2
	SeparatorTextPadding             ImVec2
	DisplayWindowPadding             ImVec2
	DisplaySafeAreaPadding           ImVec2
	DockingSeparatorSize             f32
	MouseCursorScale                 f32
	AntiAliasedLines                 bool
	AntiAliasedLinesUseTex           bool
	AntiAliasedFill                  bool
	CurveTessellationTol             f32
	CircleTessellationMaxError       f32
	Colors                           [58]ImVec4
	HoverStationaryDelay             f32
	HoverDelayShort                  f32
	HoverDelayNormal                 f32
	HoverFlagsForTooltipMouse        HoveredFlags
	HoverFlagsForTooltipNav          HoveredFlags
}



pub type KeyData = C.ImGuiKeyData
@[typedef]
struct C.ImGuiKeyData {
pub mut:
	Down             bool
	DownDuration     f32
	DownDurationPrev f32
	AnalogValue      f32
}



pub type ImVector_ImWchar = C.ImVector_ImWchar
@[typedef]
struct C.ImVector_ImWchar {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImWchar*/voidptr= unsafe{ nil }
}



pub type IO = C.ImGuiIO
@[typedef]
struct C.ImGuiIO {
pub mut:
	ConfigFlags                                   ConfigFlags
	BackendFlags                                  BackendFlags
	DisplaySize                                   ImVec2
	DeltaTime                                     f32
	IniSavingRate                                 f32
	IniFilename                                   /*&i8*/voidptr= unsafe{ nil }
	LogFilename                                   /*&i8*/voidptr= unsafe{ nil }
	UserData                                      voidptr = unsafe{ nil }
	Fonts                                         /*&ImFontAtlas*/voidptr= unsafe{ nil }
	FontGlobalScale                               f32
	FontAllowUserScaling                          bool
	FontDefault                                   /*&ImFont*/voidptr= unsafe{ nil }
	DisplayFramebufferScale                       ImVec2
	ConfigNavSwapGamepadButtons                   bool
	ConfigNavMoveSetMousePos                      bool
	ConfigNavCaptureKeyboard                      bool
	ConfigNavEscapeClearFocusItem                 bool
	ConfigNavEscapeClearFocusWindow               bool
	ConfigNavCursorVisibleAuto                    bool
	ConfigNavCursorVisibleAlways                  bool
	ConfigDockingNoSplit                          bool
	ConfigDockingWithShift                        bool
	ConfigDockingAlwaysTabBar                     bool
	ConfigDockingTransparentPayload               bool
	ConfigViewportsNoAutoMerge                    bool
	ConfigViewportsNoTaskBarIcon                  bool
	ConfigViewportsNoDecoration                   bool
	ConfigViewportsNoDefaultParent                bool
	MouseDrawCursor                               bool
	ConfigMacOSXBehaviors                         bool
	ConfigInputTrickleEventQueue                  bool
	ConfigInputTextCursorBlink                    bool
	ConfigInputTextEnterKeepActive                bool
	ConfigDragClickToInputText                    bool
	ConfigWindowsResizeFromEdges                  bool
	ConfigWindowsMoveFromTitleBarOnly             bool
	ConfigWindowsCopyContentsWithCtrlC            bool
	ConfigScrollbarScrollByPage                   bool
	ConfigMemoryCompactTimer                      f32
	MouseDoubleClickTime                          f32
	MouseDoubleClickMaxDist                       f32
	MouseDragThreshold                            f32
	KeyRepeatDelay                                f32
	KeyRepeatRate                                 f32
	ConfigErrorRecovery                           bool
	ConfigErrorRecoveryEnableAssert               bool
	ConfigErrorRecoveryEnableDebugLog             bool
	ConfigErrorRecoveryEnableTooltip              bool
	ConfigDebugIsDebuggerPresent                  bool
	ConfigDebugHighlightIdConflicts               bool
	ConfigDebugHighlightIdConflictsShowItemPicker bool
	ConfigDebugBeginReturnValueOnce               bool
	ConfigDebugBeginReturnValueLoop               bool
	ConfigDebugIgnoreFocusLoss                    bool
	ConfigDebugIniSettings                        bool
	BackendPlatformName                           /*&i8*/voidptr= unsafe{ nil }
	BackendRendererName                           /*&i8*/voidptr= unsafe{ nil }
	BackendPlatformUserData                       voidptr = unsafe{ nil }
	BackendRendererUserData                       voidptr = unsafe{ nil }
	BackendLanguageUserData                       voidptr = unsafe{ nil }
	WantCaptureMouse                              bool
	WantCaptureKeyboard                           bool
	WantTextInput                                 bool
	WantSetMousePos                               bool
	WantSaveIniSettings                           bool
	NavActive                                     bool
	NavVisible                                    bool
	Framerate                                     f32
	MetricsRenderVertices                         int
	MetricsRenderIndices                          int
	MetricsRenderWindows                          int
	MetricsActiveWindows                          int
	MouseDelta                                    ImVec2
	Ctx                                           /*&Context*/voidptr= unsafe{ nil }
	MousePos                                      ImVec2
	MouseDown                                     [5]bool
	MouseWheel                                    f32
	MouseWheelH                                   f32
	MouseSource                                   MouseSource
	MouseHoveredViewport                          ID
	KeyCtrl                                       bool
	KeyShift                                      bool
	KeyAlt                                        bool
	KeySuper                                      bool
	KeyMods                                       KeyChord
	KeysData                                      [155]KeyData
	WantCaptureMouseUnlessPopupClose              bool
	MousePosPrev                                  ImVec2
	MouseClickedPos                               [5]ImVec2
	MouseClickedTime                              [5]f64
	MouseClicked                                  [5]bool
	MouseDoubleClicked                            [5]bool
	MouseClickedCount                             [5]ImU16
	MouseClickedLastCount                         [5]ImU16
	MouseReleased                                 [5]bool
	MouseReleasedTime                             [5]f64
	MouseDownOwned                                [5]bool
	MouseDownOwnedUnlessPopupClose                [5]bool
	MouseWheelRequestAxisSwap                     bool
	MouseCtrlLeftAsRightClick                     bool
	MouseDownDuration                             [5]f32
	MouseDownDurationPrev                         [5]f32
	MouseDragMaxDistanceAbs                       [5]ImVec2
	MouseDragMaxDistanceSqr                       [5]f32
	PenPressure                                   f32
	AppFocusLost                                  bool
	AppAcceptingEvents                            bool
	InputQueueSurrogate                           ImWchar16
	InputQueueCharacters                          ImVector_ImWchar
}



pub type InputTextCallbackData = C.ImGuiInputTextCallbackData
@[typedef]
struct C.ImGuiInputTextCallbackData {
pub mut:
	Ctx            /*&Context*/voidptr= unsafe{ nil }
	EventFlag      InputTextFlags
	Flags          InputTextFlags
	UserData       voidptr = unsafe{ nil }
	EventChar      ImWchar
	EventKey       Key
	Buf            /*&i8*/voidptr= unsafe{ nil }
	BufTextLen     int
	BufSize        int
	BufDirty       bool
	CursorPos      int
	SelectionStart int
	SelectionEnd   int
}



pub type SizeCallbackData = C.ImGuiSizeCallbackData
@[typedef]
struct C.ImGuiSizeCallbackData {
pub mut:
	UserData    voidptr = unsafe{ nil }
	Pos         ImVec2
	CurrentSize ImVec2
	DesiredSize ImVec2
}



pub type WindowClass = C.ImGuiWindowClass
@[typedef]
struct C.ImGuiWindowClass {
pub mut:
	ClassId                    ID
	ParentViewportId           ID
	FocusRouteParentWindowId   ID
	ViewportFlagsOverrideSet   ViewportFlags
	ViewportFlagsOverrideClear ViewportFlags
	TabItemFlagsOverrideSet    TabItemFlags
	DockNodeFlagsOverrideSet   DockNodeFlags
	DockingAlwaysTabBar        bool
	DockingAllowUnclassed      bool
}



pub type Payload = C.ImGuiPayload
@[typedef]
struct C.ImGuiPayload {
pub mut:
	Data           voidptr = unsafe{ nil }
	DataSize       int
	SourceId       ID
	SourceParentId ID
	DataFrameCount int
	DataType       [33]i8
	Preview        bool
	Delivery       bool
}



pub type OnceUponAFrame = C.ImGuiOnceUponAFrame
@[typedef]
struct C.ImGuiOnceUponAFrame {
pub mut:
	RefFrame int
}



pub type TextRange = C.ImGuiTextRange
@[typedef]
struct C.ImGuiTextRange {
pub mut:

	b /*&i8*/voidptr= unsafe{ nil }
	e /*&i8*/voidptr= unsafe{ nil }
}



pub type ImVector_TextRange = C.ImVector_ImGuiTextRange
@[typedef]
struct C.ImVector_ImGuiTextRange {
pub mut:
	Size     int
	Capacity int
	Data     /*&TextRange*/voidptr= unsafe{ nil }
}



pub type ImVector_char = C.ImVector_char
@[typedef]
struct C.ImVector_char {
pub mut:
	Size     int
	Capacity int
	Data     /*&i8*/voidptr= unsafe{ nil }
}



pub type TextBuffer = C.ImGuiTextBuffer
@[typedef]
struct C.ImGuiTextBuffer {
pub mut:
	Buf ImVector_char
}



pub type StoragePair = C.ImGuiStoragePair
@[typedef]
struct C.ImGuiStoragePair {
pub mut:

	key ID
  val_i int
  val_f f32
  val_p voidptr
}



pub type ImVector_StoragePair = C.ImVector_ImGuiStoragePair
@[typedef]
struct C.ImVector_ImGuiStoragePair {
pub mut:
	Size     int
	Capacity int
	Data     /*&StoragePair*/voidptr= unsafe{ nil }
}



pub type Storage = C.ImGuiStorage
@[typedef]
struct C.ImGuiStorage {
pub mut:
	Data ImVector_StoragePair
}



pub type ListClipper = C.ImGuiListClipper
@[typedef]
struct C.ImGuiListClipper {
pub mut:
	Ctx              /*&Context*/voidptr= unsafe{ nil }
	DisplayStart     int
	DisplayEnd       int
	ItemsCount       int
	ItemsHeight      f32
	StartPosY        f32
	StartSeekOffsetY f64
	TempData         voidptr = unsafe{ nil }
}



pub type ImColor = C.ImColor
@[typedef]
struct C.ImColor {
pub mut:
	Value ImVec4
}

enum MultiSelectFlags_ {
 none                      = 0
 single_select             = 1 << 0
 no_select_all             = 1 << 1
 no_range_select           = 1 << 2
 no_auto_select            = 1 << 3
 no_auto_clear             = 1 << 4
 no_auto_clear_on_reselect = 1 << 5
 box_select1d              = 1 << 6
 box_select2d              = 1 << 7
 box_select_no_scroll      = 1 << 8
 clear_on_escape           = 1 << 9
 clear_on_click_void       = 1 << 10
 scope_window              = 1 << 11
 scope_rect                = 1 << 12
 select_on_click           = 1 << 13
 select_on_click_release   = 1 << 14
 nav_wrap_x                = 1 << 16
}



pub type ImVector_SelectionRequest = C.ImVector_ImGuiSelectionRequest
@[typedef]
struct C.ImVector_ImGuiSelectionRequest {
pub mut:
	Size     int
	Capacity int
	Data     /*&SelectionRequest*/voidptr= unsafe{ nil }
}



pub type MultiSelectIO = C.ImGuiMultiSelectIO
@[typedef]
struct C.ImGuiMultiSelectIO {
pub mut:
	Requests      ImVector_SelectionRequest
	RangeSrcItem  SelectionUserData
	NavIdItem     SelectionUserData
	NavIdSelected bool
	RangeSrcReset bool
	ItemsCount    int
}

enum SelectionRequestType {
 none = 0
 set_all
 set_range
}



pub type SelectionRequest = C.ImGuiSelectionRequest
@[typedef]
struct C.ImGuiSelectionRequest {
pub mut:
	Type           SelectionRequestType
	Selected       bool
	RangeDirection ImS8
	RangeFirstItem SelectionUserData
	RangeLastItem  SelectionUserData
}



pub type SelectionBasicStorage = C.ImGuiSelectionBasicStorage
@[typedef]
struct C.ImGuiSelectionBasicStorage {
pub mut:
	Size                    int
	PreserveOrder           bool
	UserData                voidptr = unsafe{ nil }
	AdapterIndexToStorageId fn (&SelectionBasicStorage, int) ID
	_SelectionOrder         int
	_Storage                Storage
}



pub type SelectionExternalStorage = C.ImGuiSelectionExternalStorage
@[typedef]
struct C.ImGuiSelectionExternalStorage {
pub mut:
	UserData               voidptr = unsafe{ nil }
	AdapterSetItemSelected fn (&SelectionExternalStorage, int, bool)
}

type ImDrawIdx = u16
type ImDrawCallback = fn (&ImDrawList, &ImDrawCmd)



pub type ImDrawCmd = C.ImDrawCmd
@[typedef]
struct C.ImDrawCmd {
pub mut:
	ClipRect               ImVec4
	TextureId              ImTextureID
	VtxOffset              u32
	IdxOffset              u32
	ElemCount              u32
	UserCallback           /*ImDrawCallback*/voidptr = unsafe{ nil }
	UserCallbackData       voidptr = unsafe{ nil }
	UserCallbackDataSize   int
	UserCallbackDataOffset int
}



pub type ImDrawVert = C.ImDrawVert
@[typedef]
struct C.ImDrawVert {
pub mut:

	pos ImVec2
	uv  ImVec2
	col ImU32
}



pub type ImDrawCmdHeader = C.ImDrawCmdHeader
@[typedef]
struct C.ImDrawCmdHeader {
pub mut:
	ClipRect  ImVec4
	TextureId ImTextureID
	VtxOffset u32
}



pub type ImVector_ImDrawCmd = C.ImVector_ImDrawCmd
@[typedef]
struct C.ImVector_ImDrawCmd {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImDrawCmd*/voidptr= unsafe{ nil }
}



pub type ImVector_ImDrawIdx = C.ImVector_ImDrawIdx
@[typedef]
struct C.ImVector_ImDrawIdx {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImDrawIdx*/voidptr= unsafe{ nil }
}



pub type ImDrawChannel = C.ImDrawChannel
@[typedef]
struct C.ImDrawChannel {
pub mut:
	_CmdBuffer ImVector_ImDrawCmd
	_IdxBuffer ImVector_ImDrawIdx
}



pub type ImVector_ImDrawChannel = C.ImVector_ImDrawChannel
@[typedef]
struct C.ImVector_ImDrawChannel {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImDrawChannel*/voidptr= unsafe{ nil }
}



pub type ImDrawListSplitter = C.ImDrawListSplitter
@[typedef]
struct C.ImDrawListSplitter {
pub mut:
	_Current  int
	_Count    int
	_Channels ImVector_ImDrawChannel
}

enum ImDrawFlags_ {
	none                       = 0
	closed                     = 1 << 0
	round_corners_top_left     = 1 << 4
	round_corners_top_right    = 1 << 5
	round_corners_bottom_left  = 1 << 6
	round_corners_bottom_right = 1 << 7
	round_corners_none         = 1 << 8
	round_corners_top          = 1 << 4 | 1 << 5
	round_corners_bottom       = 1 << 6 | 1 << 7
	round_corners_left         = 1 << 6 | 1 << 4
	round_corners_right        = 1 << 7 | 1 << 5
	round_corners_all          = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	//round_corners_default_     = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
	round_corners_mask_        = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8
}

enum ImDrawListFlags_ {
	none                       = 0
	anti_aliased_lines         = 1 << 0
	anti_aliased_lines_use_tex = 1 << 1
	anti_aliased_fill          = 1 << 2
	allow_vtx_offset           = 1 << 3
}



pub type ImVector_ImDrawVert = C.ImVector_ImDrawVert
@[typedef]
struct C.ImVector_ImDrawVert {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImDrawVert*/voidptr= unsafe{ nil }
}



pub type ImVector_ImVec2 = C.ImVector_ImVec2
@[typedef]
struct C.ImVector_ImVec2 {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImVec2*/voidptr= unsafe{ nil }
}



pub type ImVector_ImVec4 = C.ImVector_ImVec4
@[typedef]
struct C.ImVector_ImVec4 {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImVec4*/voidptr= unsafe{ nil }
}



pub type ImVector_ImTextureID = C.ImVector_ImTextureID
@[typedef]
struct C.ImVector_ImTextureID {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImTextureID*/voidptr= unsafe{ nil }
}



pub type ImVector_ImU8 = C.ImVector_ImU8
@[typedef]
struct C.ImVector_ImU8 {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImU8*/voidptr= unsafe{ nil }
}



pub type ImDrawList = C.ImDrawList
@[typedef]
struct C.ImDrawList {
pub mut:
	CmdBuffer         ImVector_ImDrawCmd
	IdxBuffer         ImVector_ImDrawIdx
	VtxBuffer         ImVector_ImDrawVert
	Flags             ImDrawListFlags
	_VtxCurrentIdx    u32
	_Data             /*&ImDrawListSharedData*/voidptr= unsafe{ nil }
	_VtxWritePtr      /*&ImDrawVert*/voidptr= unsafe{ nil }
	_IdxWritePtr      /*&ImDrawIdx*/voidptr= unsafe{ nil }
	_Path             ImVector_ImVec2
	_CmdHeader        ImDrawCmdHeader
	_Splitter         ImDrawListSplitter
	_ClipRectStack    ImVector_ImVec4
	_TextureIdStack   ImVector_ImTextureID
	_CallbacksDataBuf ImVector_ImU8
	_FringeScale      f32
	_OwnerName        /*&i8*/voidptr= unsafe{ nil }
}



pub type ImVector_ImDrawListPtr = C.ImVector_ImDrawListPtr
@[typedef]
struct C.ImVector_ImDrawListPtr {
pub mut:
	Size     int
	Capacity int
	Data     /*&&ImDrawList*/voidptr= unsafe{ nil }
}



pub type ImDrawData = C.ImDrawData
@[typedef]
struct C.ImDrawData {
pub mut:
	Valid            bool
	CmdListsCount    int
	TotalIdxCount    int
	TotalVtxCount    int
	CmdLists         ImVector_ImDrawListPtr
	DisplayPos       ImVec2
	DisplaySize      ImVec2
	FramebufferScale ImVec2
	OwnerViewport    /*&Viewport*/voidptr= unsafe{ nil }
}



pub type ImFontConfig = C.ImFontConfig
@[typedef]
struct C.ImFontConfig {
pub mut:
	FontData             voidptr = unsafe{ nil }
	FontDataSize         int
	FontDataOwnedByAtlas bool
	MergeMode            bool
	PixelSnapH           bool
	FontNo               int
	OversampleH          int
	OversampleV          int
	SizePixels           f32
	GlyphOffset          ImVec2
	GlyphRanges          /*&ImWchar*/voidptr= unsafe{ nil }
	GlyphMinAdvanceX     f32
	GlyphMaxAdvanceX     f32
	GlyphExtraAdvanceX   f32
	FontBuilderFlags     u32
	RasterizerMultiply   f32
	RasterizerDensity    f32
	EllipsisChar         ImWchar
	Name                 [40]i8
	DstFont              /*&ImFont*/voidptr= unsafe{ nil }
}



pub type ImFontGlyph = C.ImFontGlyph
@[typedef]
struct C.ImFontGlyph {
pub mut:
	Colored   u32
	Visible   u32
	Codepoint u32
	AdvanceX  f32
	X0        f32
	Y0        f32
	X1        f32
	Y1        f32
	U0        f32
	V0        f32
	U1        f32
	V1        f32
}



pub type ImVector_ImU32 = C.ImVector_ImU32
@[typedef]
struct C.ImVector_ImU32 {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImU32*/voidptr= unsafe{ nil }
}



pub type ImFontGlyphRangesBuilder = C.ImFontGlyphRangesBuilder
@[typedef]
struct C.ImFontGlyphRangesBuilder {
pub mut:
	UsedChars ImVector_ImU32
}



pub type ImFontAtlasCustomRect = C.ImFontAtlasCustomRect
@[typedef]
struct C.ImFontAtlasCustomRect {
pub mut:
	X             u16
	Y             u16
	Width         u16
	Height        u16
	GlyphID       u32
	GlyphColored  u32
	GlyphAdvanceX f32
	GlyphOffset   ImVec2
	Font          /*&ImFont*/voidptr= unsafe{ nil }
}

enum ImFontAtlasFlags_ {
	none                   = 0
	no_power_of_two_height = 1 << 0
	no_mouse_cursors       = 1 << 1
	no_baked_lines         = 1 << 2
}



pub type ImVector_ImFontPtr = C.ImVector_ImFontPtr
@[typedef]
struct C.ImVector_ImFontPtr {
pub mut:
	Size     int
	Capacity int
	Data     /*&&ImFont*/voidptr= unsafe{ nil }
}



pub type ImVector_ImFontAtlasCustomRect = C.ImVector_ImFontAtlasCustomRect
@[typedef]
struct C.ImVector_ImFontAtlasCustomRect {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImFontAtlasCustomRect*/voidptr= unsafe{ nil }
}



pub type ImVector_ImFontConfig = C.ImVector_ImFontConfig
@[typedef]
struct C.ImVector_ImFontConfig {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImFontConfig*/voidptr= unsafe{ nil }
}



pub type ImFontAtlas = C.ImFontAtlas
@[typedef]
struct C.ImFontAtlas {
pub mut:
	Flags              ImFontAtlasFlags
	TexID              ImTextureID
	TexDesiredWidth    int
	TexGlyphPadding    int
	UserData           voidptr = unsafe{ nil }
	Locked             bool
	TexReady           bool
	TexPixelsUseColors bool
	TexPixelsAlpha8    /*&u8*/voidptr= unsafe{ nil }
	TexPixelsRGBA32    /*&u32*/voidptr= unsafe{ nil }
	TexWidth           int
	TexHeight          int
	TexUvScale         ImVec2
	TexUvWhitePixel    ImVec2
	Fonts              ImVector_ImFontPtr
	CustomRects        ImVector_ImFontAtlasCustomRect
	Sources            ImVector_ImFontConfig
	TexUvLines         [33]ImVec4
	FontBuilderIO      /*&ImFontBuilderIO*/voidptr= unsafe{ nil }
	FontBuilderFlags   u32
	PackIdMouseCursors int
	PackIdLines        int
}



pub type ImVector_float = C.ImVector_float
@[typedef]
struct C.ImVector_float {
pub mut:
	Size     int
	Capacity int
	Data     /*&f32*/voidptr= unsafe{ nil }
}



pub type ImVector_ImU16 = C.ImVector_ImU16
@[typedef]
struct C.ImVector_ImU16 {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImU16*/voidptr= unsafe{ nil }
}



pub type ImVector_ImFontGlyph = C.ImVector_ImFontGlyph
@[typedef]
struct C.ImVector_ImFontGlyph {
pub mut:
	Size     int
	Capacity int
	Data     /*&ImFontGlyph*/voidptr= unsafe{ nil }
}



pub type ImFont = C.ImFont
@[typedef]
struct C.ImFont {
pub mut:
	IndexAdvanceX       ImVector_float
	FallbackAdvanceX    f32
	FontSize            f32
	IndexLookup         ImVector_ImU16
	Glyphs              ImVector_ImFontGlyph
	FallbackGlyph       /*&ImFontGlyph*/voidptr= unsafe{ nil }
	ContainerAtlas      /*&ImFontAtlas*/voidptr= unsafe{ nil }
	Sources             /*&ImFontConfig*/voidptr= unsafe{ nil }
	SourcesCount        i16
	EllipsisCharCount   i16
	EllipsisChar        ImWchar
	FallbackChar        ImWchar
	EllipsisWidth       f32
	EllipsisCharStep    f32
	Scale               f32
	Ascent              f32
	Descent             f32
	MetricsTotalSurface int
	DirtyLookupTables   bool
	Used8kPagesMap      [1]ImU8
}

enum ViewportFlags_ {
 none                   = 0
 is_platform_window     = 1 << 0
 is_platform_monitor    = 1 << 1
 owned_by_app           = 1 << 2
 no_decoration          = 1 << 3
 no_task_bar_icon       = 1 << 4
 no_focus_on_appearing  = 1 << 5
 no_focus_on_click      = 1 << 6
 no_inputs              = 1 << 7
 no_renderer_clear      = 1 << 8
 no_auto_merge          = 1 << 9
 top_most               = 1 << 10
 can_host_other_windows = 1 << 11
 is_minimized           = 1 << 12
 is_focused             = 1 << 13
}



pub type Viewport = C.ImGuiViewport
@[typedef]
struct C.ImGuiViewport {
pub mut:
	ID                    ID
	Flags                 ViewportFlags
	Pos                   ImVec2
	Size                  ImVec2
	WorkPos               ImVec2
	WorkSize              ImVec2
	DpiScale              f32
	ParentViewportId      ID
	DrawData              /*&ImDrawData*/voidptr= unsafe{ nil }
	RendererUserData      voidptr = unsafe{ nil }
	PlatformUserData      voidptr = unsafe{ nil }
	PlatformHandle        voidptr = unsafe{ nil }
	PlatformHandleRaw     voidptr = unsafe{ nil }
	PlatformWindowCreated bool
	PlatformRequestMove   bool
	PlatformRequestResize bool
	PlatformRequestClose  bool
}



pub type ImVector_PlatformMonitor = C.ImVector_ImGuiPlatformMonitor
@[typedef]
struct C.ImVector_ImGuiPlatformMonitor {
pub mut:
	Size     int
	Capacity int
	Data     /*&PlatformMonitor*/voidptr= unsafe{ nil }
}



pub type ImVector_ViewportPtr = C.ImVector_ImGuiViewportPtr
@[typedef]
struct C.ImVector_ImGuiViewportPtr {
pub mut:
	Size     int
	Capacity int
	Data     /*&&Viewport*/voidptr= unsafe{ nil }
}



pub type PlatformIO = C.ImGuiPlatformIO
@[typedef]
struct C.ImGuiPlatformIO {
pub mut:
	Platform_GetClipboardTextFn      fn (&Context) &i8
	Platform_SetClipboardTextFn      fn (&Context, &i8)
	Platform_ClipboardUserData       voidptr = unsafe{ nil }
	Platform_OpenInShellFn           fn (&Context, &i8) bool
	Platform_OpenInShellUserData     voidptr = unsafe{ nil }
	Platform_SetImeDataFn            fn (&Context, &Viewport, &PlatformImeData)
	Platform_ImeUserData             voidptr = unsafe{ nil }
	Platform_LocaleDecimalPoint      ImWchar
	Renderer_RenderState             voidptr = unsafe{ nil }
	Platform_CreateWindow            fn (&Viewport)
	Platform_DestroyWindow           fn (&Viewport)
	Platform_ShowWindow              fn (&Viewport)
	Platform_SetWindowPos            fn (&Viewport, ImVec2)
	Platform_GetWindowPos            fn (&Viewport) ImVec2
	Platform_SetWindowSize           fn (&Viewport, ImVec2)
	Platform_GetWindowSize           fn (&Viewport) ImVec2
	Platform_SetWindowFocus          fn (&Viewport)
	Platform_GetWindowFocus          fn (&Viewport) bool
	Platform_GetWindowMinimized      fn (&Viewport) bool
	Platform_SetWindowTitle          fn (&Viewport, &i8)
	Platform_SetWindowAlpha          fn (&Viewport, f32)
	Platform_UpdateWindow            fn (&Viewport)
	Platform_RenderWindow            fn (&Viewport, voidptr)
	Platform_SwapBuffers             fn (&Viewport, voidptr)
	Platform_GetWindowDpiScale       fn (&Viewport) f32
	Platform_OnChangedViewport       fn (&Viewport)
	Platform_GetWindowWorkAreaInsets fn (&Viewport) ImVec4
	Platform_CreateVkSurface         fn (&Viewport, ImU64, voidptr, &ImU64) int
	Renderer_CreateWindow            fn (&Viewport)
	Renderer_DestroyWindow           fn (&Viewport)
	Renderer_SetWindowSize           fn (&Viewport, ImVec2)
	Renderer_RenderWindow            fn (&Viewport, voidptr)
	Renderer_SwapBuffers             fn (&Viewport, voidptr)
	Monitors                         ImVector_PlatformMonitor
	Viewports                        ImVector_ViewportPtr
}



pub type PlatformMonitor = C.ImGuiPlatformMonitor
@[typedef]
struct C.ImGuiPlatformMonitor {
pub mut:
	MainPos        ImVec2
	MainSize       ImVec2
	WorkPos        ImVec2
	WorkSize       ImVec2
	DpiScale       f32
	PlatformHandle voidptr = unsafe{ nil }
}



pub type PlatformImeData = C.ImGuiPlatformImeData
@[typedef]
struct C.ImGuiPlatformImeData {
pub mut:
	WantVisible     bool
	InputPos        ImVec2
	InputLineHeight f32
}

type DataAuthority = int
type LayoutType = int
type ActivateFlags = int
type DebugLogFlags = int
type FocusRequestFlags = int
type ItemStatusFlags = int
type OldColumnFlags = int
type LogFlags = int
type NavRenderCursorFlags = int
type NavMoveFlags = int
type NextItemDataFlags = int
type NextWindowDataFlags = int
type ScrollFlags = int
type SeparatorFlags = int
type TextFlags = int
type TooltipFlags = int
type TypingSelectFlags = int
type WindowRefreshFlags = int

/*
@[weak]
__global G &Context
*/
pub type ImFileHandle = &voidptr



pub type ImVec1 = C.ImVec1
@[typedef]
struct C.ImVec1 {
pub mut:

	x f32
}



pub type ImVec2ih = C.ImVec2ih
@[typedef]
struct C.ImVec2ih {
pub mut:

	x i16
	y i16
}



pub type ImRect = C.ImRect
@[typedef]
struct C.ImRect {
pub mut:
	Min ImVec2
	Max ImVec2
}

type ImBitArrayPtr = &u32



pub type ImBitVector = C.ImBitVector
@[typedef]
struct C.ImBitVector {
pub mut:
	Storage ImVector_ImU32
}

type ImPoolIdx = int



pub type ImVector_int = C.ImVector_int
@[typedef]
struct C.ImVector_int {
pub mut:
	Size     int
	Capacity int
	Data     /*&int*/voidptr= unsafe{ nil }
}



pub type TextIndex = C.ImGuiTextIndex
@[typedef]
struct C.ImGuiTextIndex {
pub mut:
	LineOffsets ImVector_int
	EndOffset   int
}



pub type ImDrawListSharedData = C.ImDrawListSharedData
@[typedef]
struct C.ImDrawListSharedData {
pub mut:
	TexUvWhitePixel       ImVec2
	TexUvLines            /*&ImVec4*/voidptr= unsafe{ nil }
	Font                  /*&ImFont*/voidptr= unsafe{ nil }
	FontSize              f32
	FontScale             f32
	CurveTessellationTol  f32
	CircleSegmentMaxError f32
	InitialFringeScale    f32
	InitialFlags          ImDrawListFlags
	ClipRectFullscreen    ImVec4
	TempBuffer            ImVector_ImVec2
	ArcFastVtx            [48]ImVec2
	ArcFastRadiusCutoff   f32
	CircleSegmentCounts   [64]ImU8
}



pub type ImDrawDataBuilder = C.ImDrawDataBuilder
@[typedef]
struct C.ImDrawDataBuilder {
pub mut:
	Layers     [2]&ImVector_ImDrawListPtr
	LayerData1 ImVector_ImDrawListPtr
}



pub type StyleVarInfo = C.ImGuiStyleVarInfo
@[typedef]
struct C.ImGuiStyleVarInfo {
pub mut:
	Count    ImU32
	DataType DataType
	Offset   ImU32
}



pub type ColorMod = C.ImGuiColorMod
@[typedef]
struct C.ImGuiColorMod {
pub mut:
	Col         Col
	BackupValue ImVec4
}



pub type StyleMod = C.ImGuiStyleMod
@[typedef]
struct C.ImGuiStyleMod {
pub mut:
	VarIdx StyleVar
  BackupInt [2]int
  BackupFloat [2]f32
}



pub type DataTypeStorage = C.ImGuiDataTypeStorage
@[typedef]
struct C.ImGuiDataTypeStorage {
pub mut:
	Data [8]ImU8
}



pub type DataTypeInfo = C.ImGuiDataTypeInfo
@[typedef]
struct C.ImGuiDataTypeInfo {
pub mut:
	Size     usize
	Name     /*&i8*/voidptr= unsafe{ nil }
	PrintFmt /*&i8*/voidptr= unsafe{ nil }
	ScanFmt  /*&i8*/voidptr= unsafe{ nil }
}

enum DataTypePrivate_ {
 pointer = int(DataType_.count)
 id
}

enum ItemFlagsPrivate_ {
 disabled                   = 1 << 10
 read_only                  = 1 << 11
 mixed_value                = 1 << 12
 no_window_hoverable_check  = 1 << 13
 allow_overlap              = 1 << 14
 no_nav_disable_mouse_hover = 1 << 15
 no_mark_edited             = 1 << 16
 inputable                  = 1 << 20
 has_selection_user_data    = 1 << 21
 is_multi_select            = 1 << 22
 default_                   = 1 << 4
}

enum ItemStatusFlags_ {
 none              = 0
 hovered_rect      = 1 << 0
 has_display_rect  = 1 << 1
 edited            = 1 << 2
 toggled_selection = 1 << 3
 toggled_open      = 1 << 4
 has_deactivated   = 1 << 5
 deactivated       = 1 << 6
 hovered_window    = 1 << 7
 visible           = 1 << 8
 has_clip_rect     = 1 << 9
 has_shortcut      = 1 << 10
}

enum HoveredFlagsPrivate_ {
 delay_mask_                        = 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
 allowed_mask_for_is_window_hovered = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 7 | 1 << 12 | 1 << 13
 allowed_mask_for_is_item_hovered   = 1 << 5 | 1 << 7 | 1 << 8 | 1 << 9 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
}

enum InputTextFlagsPrivate_ {
 multiline              = 1 << 26
 merged_item            = 1 << 27
 localize_decimal_point = 1 << 28
}

enum ButtonFlagsPrivate_ {
 pressed_on_click                  = 1 << 4
 pressed_on_click_release          = 1 << 5
 pressed_on_click_release_anywhere = 1 << 6
 pressed_on_release                = 1 << 7
 pressed_on_double_click           = 1 << 8
 pressed_on_drag_drop_hold         = 1 << 9
 flatten_children                  = 1 << 11
 allow_overlap                     = 1 << 12
 align_text_base_line              = 1 << 15
 no_key_mods_allowed               = 1 << 16
 no_holding_active_id              = 1 << 17
 no_nav_focus                      = 1 << 18
 no_hovered_on_focus               = 1 << 19
 no_set_key_owner                  = 1 << 20
 no_test_key_owner                 = 1 << 21
 pressed_on_mask_                  = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8 | 1 << 9
 //pressed_on_default_               = 1 << 5
}

enum ComboFlagsPrivate_ {
 custom_preview = 1 << 20
}

enum SliderFlagsPrivate_ {
 vertical  = 1 << 20
 read_only = 1 << 21
}

enum SelectableFlagsPrivate_ {
 no_holding_active_id     = 1 << 20
 select_on_nav            = 1 << 21
 select_on_click          = 1 << 22
 select_on_release        = 1 << 23
 span_avail_width         = 1 << 24
 set_nav_id_on_hover      = 1 << 25
 no_pad_with_half_spacing = 1 << 26
 no_set_key_owner         = 1 << 27
}

enum TreeNodeFlagsPrivate_ {
 clip_label_for_trailing_button = 1 << 28
 upside_down_arrow              = 1 << 29
 open_on_mask_                  = 1 << 6 | 1 << 7
}

enum SeparatorFlags_ {
 none             = 0
 horizontal       = 1 << 0
 vertical         = 1 << 1
 span_all_columns = 1 << 2
}

enum FocusRequestFlags_ {
 none                  = 0
 restore_focused_child = 1 << 0
 unless_below_modal    = 1 << 1
}

enum TextFlags_ {
 none                            = 0
 no_width_for_large_clipped_text = 1 << 0
}

enum TooltipFlags_ {
 none              = 0
 override_previous = 1 << 1
}

enum LayoutType_ {
 horizontal = 0
 vertical   = 1
}

enum LogFlags_ {
 none             = 0
 output_tty       = 1 << 0
 output_file      = 1 << 1
 output_buffer    = 1 << 2
 output_clipboard = 1 << 3
 output_mask_     = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
}

enum Axis {
 none = -1
 x    = 0
 y    = 1
}

enum PlotType {
 lines
 histogram
}



pub type ComboPreviewData = C.ImGuiComboPreviewData
@[typedef]
struct C.ImGuiComboPreviewData {
pub mut:
	PreviewRect                  ImRect
	BackupCursorPos              ImVec2
	BackupCursorMaxPos           ImVec2
	BackupCursorPosPrevLine      ImVec2
	BackupPrevLineTextBaseOffset f32
	BackupLayout                 LayoutType
}



pub type GroupData = C.ImGuiGroupData
@[typedef]
struct C.ImGuiGroupData {
pub mut:
	WindowID                     ID
	BackupCursorPos              ImVec2
	BackupCursorMaxPos           ImVec2
	BackupCursorPosPrevLine      ImVec2
	BackupIndent                 ImVec1
	BackupGroupOffset            ImVec1
	BackupCurrLineSize           ImVec2
	BackupCurrLineTextBaseOffset f32
	BackupActiveIdIsAlive        ID
	BackupDeactivatedIdIsAlive   bool
	BackupHoveredIdIsAlive       bool
	BackupIsSameLine             bool
	EmitItem                     bool
}



pub type MenuColumns = C.ImGuiMenuColumns
@[typedef]
struct C.ImGuiMenuColumns {
pub mut:
	TotalWidth     ImU32
	NextTotalWidth ImU32
	Spacing        ImU16
	OffsetIcon     ImU16
	OffsetLabel    ImU16
	OffsetShortcut ImU16
	OffsetMark     ImU16
	Widths         [4]ImU16
}



pub type InputTextDeactivatedState = C.ImGuiInputTextDeactivatedState
@[typedef]
struct C.ImGuiInputTextDeactivatedState {
pub mut:
	ID    ID
	TextA ImVector_char
}


pub type ImStbTexteditState = C.STB_TexteditState
@[typedef]
struct C.STB_TexteditState {}



pub type InputTextState = C.ImGuiInputTextState
@[typedef]
struct C.ImGuiInputTextState {
pub mut:
	Ctx                  /*&Context*/voidptr= unsafe{ nil }
	Stb                  /*&ImStbTexteditState*/voidptr= unsafe{ nil }
	Flags                InputTextFlags
	ID                   ID
	TextLen              int
	TextSrc              /*&i8*/voidptr= unsafe{ nil }
	TextA                ImVector_char
	TextToRevertTo       ImVector_char
	CallbackTextBackup   ImVector_char
	BufCapacity          int
	Scroll               ImVec2
	CursorAnim           f32
	CursorFollow         bool
	SelectedAllMouseLock bool
	Edited               bool
	WantReloadUserBuf    bool
	ReloadSelectionStart int
	ReloadSelectionEnd   int
}

enum WindowRefreshFlags_ {
 none                 = 0
 try_to_avoid_refresh = 1 << 0
 refresh_on_hover     = 1 << 1
 refresh_on_focus     = 1 << 2
}

enum NextWindowDataFlags_ {
 none                = 0
 has_pos             = 1 << 0
 has_size            = 1 << 1
 has_content_size    = 1 << 2
 has_collapsed       = 1 << 3
 has_size_constraint = 1 << 4
 has_focus           = 1 << 5
 has_bg_alpha        = 1 << 6
 has_scroll          = 1 << 7
 has_window_flags    = 1 << 8
 has_child_flags     = 1 << 9
 has_refresh_policy  = 1 << 10
 has_viewport        = 1 << 11
 has_dock            = 1 << 12
 has_window_class    = 1 << 13
}



pub type NextWindowData = C.ImGuiNextWindowData
@[typedef]
struct C.ImGuiNextWindowData {
pub mut:
	HasFlags             NextWindowDataFlags
	PosCond              Cond
	SizeCond             Cond
	CollapsedCond        Cond
	DockCond             Cond
	PosVal               ImVec2
	PosPivotVal          ImVec2
	SizeVal              ImVec2
	ContentSizeVal       ImVec2
	ScrollVal            ImVec2
	WindowFlags          WindowFlags
	ChildFlags           ChildFlags
	PosUndock            bool
	CollapsedVal         bool
	SizeConstraintRect   ImRect
	SizeCallback         /*SizeCallback*/voidptr = unsafe{ nil }
	SizeCallbackUserData voidptr = unsafe{ nil }
	BgAlphaVal           f32
	ViewportId           ID
	DockId               ID
	WindowClass          WindowClass
	MenuBarOffsetMinVal  ImVec2
	RefreshFlagsVal      WindowRefreshFlags
}

enum NextItemDataFlags_ {
 none           = 0
 has_width      = 1 << 0
 has_open       = 1 << 1
 has_shortcut   = 1 << 2
 has_ref_val    = 1 << 3
 has_storage_id = 1 << 4
}



pub type NextItemData = C.ImGuiNextItemData
@[typedef]
struct C.ImGuiNextItemData {
pub mut:
	HasFlags          NextItemDataFlags
	ItemFlags         ItemFlags
	FocusScopeId      ID
	SelectionUserData SelectionUserData
	Width             f32
	Shortcut          KeyChord
	ShortcutFlags     InputFlags
	OpenVal           bool
	OpenCond          ImU8
	RefVal            DataTypeStorage
	StorageId         ID
}



pub type LastItemData = C.ImGuiLastItemData
@[typedef]
struct C.ImGuiLastItemData {
pub mut:
	ID          ID
	ItemFlags   ItemFlags
	StatusFlags ItemStatusFlags
	Rect        ImRect
	NavRect     ImRect
	DisplayRect ImRect
	ClipRect    ImRect
	Shortcut    KeyChord
}



pub type TreeNodeStackData = C.ImGuiTreeNodeStackData
@[typedef]
struct C.ImGuiTreeNodeStackData {
pub mut:
	ID        ID
	TreeFlags TreeNodeFlags
	ItemFlags ItemFlags
	NavRect   ImRect
}



pub type ErrorRecoveryState = C.ImGuiErrorRecoveryState
@[typedef]
struct C.ImGuiErrorRecoveryState {
pub mut:
	SizeOfWindowStack     i16
	SizeOfIDStack         i16
	SizeOfTreeStack       i16
	SizeOfColorStack      i16
	SizeOfStyleVarStack   i16
	SizeOfFontStack       i16
	SizeOfFocusScopeStack i16
	SizeOfGroupStack      i16
	SizeOfItemFlagsStack  i16
	SizeOfBeginPopupStack i16
	SizeOfDisabledStack   i16
}



pub type WindowStackData = C.ImGuiWindowStackData
@[typedef]
struct C.ImGuiWindowStackData {
pub mut:
	Window                              /*&Window*/voidptr= unsafe{ nil }
	ParentLastItemDataBackup            LastItemData
	StackSizesInBegin                   ErrorRecoveryState
	DisabledOverrideReenable            bool
	DisabledOverrideReenableAlphaBackup f32
}



pub type ShrinkWidthItem = C.ImGuiShrinkWidthItem
@[typedef]
struct C.ImGuiShrinkWidthItem {
pub mut:
	Index        int
	Width        f32
	InitialWidth f32
}



pub type PtrOrIndex = C.ImGuiPtrOrIndex
@[typedef]
struct C.ImGuiPtrOrIndex {
pub mut:
	Ptr   voidptr = unsafe{ nil }
	Index int
}



pub type DeactivatedItemData = C.ImGuiDeactivatedItemData
@[typedef]
struct C.ImGuiDeactivatedItemData {
pub mut:
	ID                  ID
	ElapseFrame         int
	HasBeenEditedBefore bool
	IsAlive             bool
}

enum PopupPositionPolicy {
 default
 combo_box
 tooltip
}



pub type PopupData = C.ImGuiPopupData
@[typedef]
struct C.ImGuiPopupData {
pub mut:
	PopupId          ID
	Window           /*&Window*/voidptr= unsafe{ nil }
	RestoreNavWindow /*&Window*/voidptr= unsafe{ nil }
	ParentNavLayer   int
	OpenFrameCount   int
	OpenParentId     ID
	OpenPopupPos     ImVec2
	OpenMousePos     ImVec2
}



pub type ImBitArray_Key_NamedKey_COUNT__lessKey_NamedKey_BEGIN = C.ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN
@[typedef]
struct C.ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN {
pub mut:
	Storage [5]ImU32
}

type ImBitArrayForNamedKeys = C.ImBitArray_ImGuiKey_NamedKey_COUNT__lessImGuiKey_NamedKey_BEGIN

enum InputEventType {
 none = 0
 mouse_pos
 mouse_wheel
 mouse_button
 mouse_viewport
 key
 text
 focus
 count
}

enum InputSource {
 none = 0
 mouse
 keyboard
 gamepad
 count
}



pub type InputEventMousePos = C.ImGuiInputEventMousePos
@[typedef]
struct C.ImGuiInputEventMousePos {
pub mut:
	PosX        f32
	PosY        f32
	MouseSource MouseSource
}



pub type InputEventMouseWheel = C.ImGuiInputEventMouseWheel
@[typedef]
struct C.ImGuiInputEventMouseWheel {
pub mut:
	WheelX      f32
	WheelY      f32
	MouseSource MouseSource
}



pub type InputEventMouseButton = C.ImGuiInputEventMouseButton
@[typedef]
struct C.ImGuiInputEventMouseButton {
pub mut:
	Button      int
	Down        bool
	MouseSource MouseSource
}



pub type InputEventMouseViewport = C.ImGuiInputEventMouseViewport
@[typedef]
struct C.ImGuiInputEventMouseViewport {
pub mut:
	HoveredViewportID ID
}



pub type InputEventKey = C.ImGuiInputEventKey
@[typedef]
struct C.ImGuiInputEventKey {
pub mut:
	Key         Key
	Down        bool
	AnalogValue f32
}



pub type InputEventText = C.ImGuiInputEventText
@[typedef]
struct C.ImGuiInputEventText {
pub mut:
	Char u32
}



pub type InputEventAppFocused = C.ImGuiInputEventAppFocused
@[typedef]
struct C.ImGuiInputEventAppFocused {
pub mut:
	Focused bool
}



pub type InputEvent = C.ImGuiInputEvent
@[typedef]
struct C.ImGuiInputEvent {
pub mut:
	Type              InputEventType
	Source            InputSource
	EventId           ImU32
	AddedByTestEngine bool
}

type KeyRoutingIndex = i16



pub type KeyRoutingData = C.ImGuiKeyRoutingData
@[typedef]
struct C.ImGuiKeyRoutingData {
pub mut:
	NextEntryIndex   KeyRoutingIndex
	Mods             ImU16
	RoutingCurrScore ImU8
	RoutingNextScore ImU8
	RoutingCurr      ID
	RoutingNext      ID
}



pub type ImVector_KeyRoutingData = C.ImVector_ImGuiKeyRoutingData
@[typedef]
struct C.ImVector_ImGuiKeyRoutingData {
pub mut:
	Size     int
	Capacity int
	Data     /*&KeyRoutingData*/voidptr= unsafe{ nil }
}



pub type KeyRoutingTable = C.ImGuiKeyRoutingTable
@[typedef]
struct C.ImGuiKeyRoutingTable {
pub mut:
	Index       [155]KeyRoutingIndex
	Entries     ImVector_KeyRoutingData
	EntriesNext ImVector_KeyRoutingData
}



pub type KeyOwnerData = C.ImGuiKeyOwnerData
@[typedef]
struct C.ImGuiKeyOwnerData {
pub mut:
	OwnerCurr        ID
	OwnerNext        ID
	LockThisFrame    bool
	LockUntilRelease bool
}

enum InputFlagsPrivate_ {
 repeat_rate_default                    = 1 << 1
 repeat_rate_nav_move                   = 1 << 2
 repeat_rate_nav_tweak                  = 1 << 3
 repeat_until_release                   = 1 << 4
 repeat_until_key_mods_change           = 1 << 5
 repeat_until_key_mods_change_from_none = 1 << 6
 repeat_until_other_key_press           = 1 << 7
 lock_this_frame                        = 1 << 20
 lock_until_release                     = 1 << 21
 cond_hovered                           = 1 << 22
 cond_active                            = 1 << 23
 /* cond_default_                          = 1 << 22 | cond_active */
 repeat_rate_mask_                      = 1 << 1 | 1 << 2 | 1 << 3
 repeat_until_mask_                     = 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
 repeat_mask_                           = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7
 cond_mask_                             = 1 << 22 | 1 << 23
 route_type_mask_                       = 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13
 route_options_mask_                    = 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
 /* supported_by_is_key_pressed            = repeat_mask_ */
 supported_by_is_mouse_clicked          = 1 << 0
 supported_by_shortcut                  = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17
 supported_by_set_next_item_shortcut    = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15 | 1 << 16 | 1 << 17 | 1 << 18
 supported_by_set_key_owner             = 1 << 20 | 1 << 21
 supported_by_set_item_key_owner        = 1 << 20 | 1 << 21 | 1 << 22 | 1 << 23
}



pub type ListClipperRange = C.ImGuiListClipperRange
@[typedef]
struct C.ImGuiListClipperRange {
pub mut:
	Min                 int
	Max                 int
	PosToIndexConvert   bool
	PosToIndexOffsetMin ImS8
	PosToIndexOffsetMax ImS8
}



pub type ImVector_ListClipperRange = C.ImVector_ImGuiListClipperRange
@[typedef]
struct C.ImVector_ImGuiListClipperRange {
pub mut:
	Size     int
	Capacity int
	Data     /*&ListClipperRange*/voidptr= unsafe{ nil }
}



pub type ListClipperData = C.ImGuiListClipperData
@[typedef]
struct C.ImGuiListClipperData {
pub mut:
	ListClipper     /*&ListClipper*/voidptr= unsafe{ nil }
	LossynessOffset f32
	StepNo          int
	ItemsFrozen     int
	Ranges          ImVector_ListClipperRange
}

enum ActivateFlags_ {
 none                  = 0
 prefer_input          = 1 << 0
 prefer_tweak          = 1 << 1
 try_to_preserve_state = 1 << 2
 from_tabbing          = 1 << 3
 from_shortcut         = 1 << 4
}

enum ScrollFlags_ {
 none                  = 0
 keep_visible_edge_x   = 1 << 0
 keep_visible_edge_y   = 1 << 1
 keep_visible_center_x = 1 << 2
 keep_visible_center_y = 1 << 3
 always_center_x       = 1 << 4
 always_center_y       = 1 << 5
 no_scroll_parent      = 1 << 6
 mask_x_               = 1 << 0 | 1 << 2 | 1 << 4
 mask_y_               = 1 << 1 | 1 << 3 | 1 << 5
}

enum NavRenderCursorFlags_ {
 none        = 0
 compact     = 1 << 1
 always_draw = 1 << 2
 no_rounding = 1 << 3
}

enum NavMoveFlags_ {
 none                      = 0
 loop_x                    = 1 << 0
 loop_y                    = 1 << 1
 wrap_x                    = 1 << 2
 wrap_y                    = 1 << 3
 wrap_mask_                = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3
 allow_current_nav_id      = 1 << 4
 also_score_visible_set    = 1 << 5
 scroll_to_edge_y          = 1 << 6
 forwarded                 = 1 << 7
 debug_no_result           = 1 << 8
 focus_api                 = 1 << 9
 is_tabbing                = 1 << 10
 is_page_move              = 1 << 11
 activate                  = 1 << 12
 no_select                 = 1 << 13
 no_set_nav_cursor_visible = 1 << 14
 no_clear_active_id        = 1 << 15
}

enum NavLayer {
 main = 0
 menu = 1
 count
}



pub type NavItemData = C.ImGuiNavItemData
@[typedef]
struct C.ImGuiNavItemData {
pub mut:
	Window            /*&Window*/voidptr= unsafe{ nil }
	ID                ID
	FocusScopeId      ID
	RectRel           ImRect
	ItemFlags         ItemFlags
	DistBox           f32
	DistCenter        f32
	DistAxial         f32
	SelectionUserData SelectionUserData
}



pub type FocusScopeData = C.ImGuiFocusScopeData
@[typedef]
struct C.ImGuiFocusScopeData {
pub mut:
	ID       ID
	WindowID ID
}

enum TypingSelectFlags_ {
 none                   = 0
 allow_backspace        = 1 << 0
 allow_single_char_mode = 1 << 1
}



pub type TypingSelectRequest = C.ImGuiTypingSelectRequest
@[typedef]
struct C.ImGuiTypingSelectRequest {
pub mut:
	Flags           TypingSelectFlags
	SearchBufferLen int
	SearchBuffer    /*&i8*/voidptr= unsafe{ nil }
	SelectRequest   bool
	SingleCharMode  bool
	SingleCharSize  ImS8
}



pub type TypingSelectState = C.ImGuiTypingSelectState
@[typedef]
struct C.ImGuiTypingSelectState {
pub mut:
	Request            TypingSelectRequest
	SearchBuffer       [64]i8
	FocusScope         ID
	LastRequestFrame   int
	LastRequestTime    f32
	SingleCharModeLock bool
}

enum OldColumnFlags_ {
 none                      = 0
 no_border                 = 1 << 0
 no_resize                 = 1 << 1
 no_preserve_widths        = 1 << 2
 no_force_within_window    = 1 << 3
 grow_parent_contents_size = 1 << 4
}



pub type OldColumnData = C.ImGuiOldColumnData
@[typedef]
struct C.ImGuiOldColumnData {
pub mut:
	OffsetNorm             f32
	OffsetNormBeforeResize f32
	Flags                  OldColumnFlags
	ClipRect               ImRect
}



pub type ImVector_OldColumnData = C.ImVector_ImGuiOldColumnData
@[typedef]
struct C.ImVector_ImGuiOldColumnData {
pub mut:
	Size     int
	Capacity int
	Data     /*&OldColumnData*/voidptr= unsafe{ nil }
}



pub type OldColumns = C.ImGuiOldColumns
@[typedef]
struct C.ImGuiOldColumns {
pub mut:
	ID                       ID
	Flags                    OldColumnFlags
	IsFirstFrame             bool
	IsBeingResized           bool
	Current                  int
	Count                    int
	OffMinX                  f32
	OffMaxX                  f32
	LineMinY                 f32
	LineMaxY                 f32
	HostCursorPosY           f32
	HostCursorMaxPosX        f32
	HostInitialClipRect      ImRect
	HostBackupClipRect       ImRect
	HostBackupParentWorkRect ImRect
	Columns                  ImVector_OldColumnData
	Splitter                 ImDrawListSplitter
}



pub type BoxSelectState = C.ImGuiBoxSelectState
@[typedef]
struct C.ImGuiBoxSelectState {
pub mut:
	ID                    ID
	IsActive              bool
	IsStarting            bool
	IsStartedFromVoid     bool
	IsStartedSetNavIdOnce bool
	RequestClear          bool
	KeyMods               KeyChord
	StartPosRel           ImVec2
	EndPosRel             ImVec2
	ScrollAccum           ImVec2
	Window                /*&Window*/voidptr= unsafe{ nil }
	UnclipMode            bool
	UnclipRect            ImRect
	BoxSelectRectPrev     ImRect
	BoxSelectRectCurr     ImRect
}



pub type MultiSelectTempData = C.ImGuiMultiSelectTempData
@[typedef]
struct C.ImGuiMultiSelectTempData {
pub mut:
	IO                 MultiSelectIO
	Storage            /*&MultiSelectState*/voidptr= unsafe{ nil }
	FocusScopeId       ID
	Flags              MultiSelectFlags
	ScopeRectMin       ImVec2
	BackupCursorMaxPos ImVec2
	LastSubmittedItem  SelectionUserData
	BoxSelectId        ID
	KeyMods            KeyChord
	LoopRequestSetAll  ImS8
	IsEndIO            bool
	IsFocused          bool
	IsKeyboardSetRange bool
	NavIdPassedBy      bool
	RangeSrcPassedBy   bool
	RangeDstPassedBy   bool
}



pub type MultiSelectState = C.ImGuiMultiSelectState
@[typedef]
struct C.ImGuiMultiSelectState {
pub mut:
	Window            /*&Window*/voidptr= unsafe{ nil }
	ID                ID
	LastFrameActive   int
	LastSelectionSize int
	RangeSelected     ImS8
	NavIdSelected     ImS8
	RangeSrcItem      SelectionUserData
	NavIdItem         SelectionUserData
}

enum DockNodeFlagsPrivate_ {
 dock_space                    = 1 << 10
 central_node                  = 1 << 11
 no_tab_bar                    = 1 << 12
 hidden_tab_bar                = 1 << 13
 no_window_menu_button         = 1 << 14
 no_close_button               = 1 << 15
 no_resize_x                   = 1 << 16
 no_resize_y                   = 1 << 17
 docked_windows_in_focus_route = 1 << 18
 no_docking_split_other        = 1 << 19
 no_docking_over_me            = 1 << 20
 no_docking_over_other         = 1 << 21
 no_docking_over_empty         = 1 << 22
 no_docking                    = 1 << 20 | 1 << 21 | 1 << 22 | 1 << 4 | 1 << 19
 shared_flags_inherit_mask_    = int(~0)
 no_resize_flags_mask_         = 1 << 5 | 1 << 16 | 1 << 17
 local_flags_transfer_mask_    = 1 << 4 | 1 << 5 | 1 << 16 | 1 << 17 | 1 << 6 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15
 saved_flags_mask_             = 1 << 5 | 1 << 16 | 1 << 17 | 1 << 10 | 1 << 11 | 1 << 12 | 1 << 13 | 1 << 14 | 1 << 15
}

enum DataAuthority_ {
 auto
 dock_node
 window
}

enum DockNodeState {
 unknown
 host_window_hidden_because_single_window
 host_window_hidden_because_windows_are_resizing
 host_window_visible
}



pub type ImVector_WindowPtr = C.ImVector_ImGuiWindowPtr
@[typedef]
struct C.ImVector_ImGuiWindowPtr {
pub mut:
	Size     int
	Capacity int
	Data     /*&&Window*/voidptr= unsafe{ nil }
}



pub type DockNode = C.ImGuiDockNode
@[typedef]
struct C.ImGuiDockNode {
pub mut:
	ID                     ID
	SharedFlags            DockNodeFlags
	LocalFlags             DockNodeFlags
	LocalFlagsInWindows    DockNodeFlags
	MergedFlags            DockNodeFlags
	State                  DockNodeState
	ParentNode             /*&DockNode*/voidptr= unsafe{ nil }
	ChildNodes             [2]&DockNode
	Windows                ImVector_WindowPtr
	TabBar                 /*&TabBar*/voidptr= unsafe{ nil }
	Pos                    ImVec2
	Size                   ImVec2
	SizeRef                ImVec2
	SplitAxis              Axis
	WindowClass            WindowClass
	LastBgColor            ImU32
	HostWindow             /*&Window*/voidptr= unsafe{ nil }
	VisibleWindow          /*&Window*/voidptr= unsafe{ nil }
	CentralNode            /*&DockNode*/voidptr= unsafe{ nil }
	OnlyNodeWithWindows    /*&DockNode*/voidptr= unsafe{ nil }
	CountNodeWithWindows   int
	LastFrameAlive         int
	LastFrameActive        int
	LastFrameFocused       int
	LastFocusedNodeId      ID
	SelectedTabId          ID
	WantCloseTabId         ID
	RefViewportId          ID
	AuthorityForPos        DataAuthority
	AuthorityForSize       DataAuthority
	AuthorityForViewport   DataAuthority
	IsVisible              bool
	IsFocused              bool
	IsBgDrawnThisFrame     bool
	HasCloseButton         bool
	HasWindowMenuButton    bool
	HasCentralNodeChild    bool
	WantCloseAll           bool
	WantLockSizeOnce       bool
	WantMouseMove          bool
	WantHiddenTabBarUpdate bool
	WantHiddenTabBarToggle bool
}

enum WindowDockStyleCol {
 text
 tab_hovered
 tab_focused
 tab_selected
 tab_selected_overline
 tab_dimmed
 tab_dimmed_selected
 tab_dimmed_selected_overline
 count
}



pub type WindowDockStyle = C.ImGuiWindowDockStyle
@[typedef]
struct C.ImGuiWindowDockStyle {
pub mut:
	Colors [8]ImU32
}



pub type ImVector_DockRequest = C.ImVector_ImGuiDockRequest
@[typedef]
struct C.ImVector_ImGuiDockRequest {
pub mut:
	Size     int
	Capacity int
	Data     /*&DockRequest*/voidptr= unsafe{ nil }
}



pub type ImVector_DockNodeSettings = C.ImVector_ImGuiDockNodeSettings
@[typedef]
struct C.ImVector_ImGuiDockNodeSettings {
pub mut:
	Size     int
	Capacity int
	Data     /*&DockNodeSettings*/voidptr= unsafe{ nil }
}



pub type DockContext = C.ImGuiDockContext
@[typedef]
struct C.ImGuiDockContext {
pub mut:
	Nodes           Storage
	Requests        ImVector_DockRequest
	NodesSettings   ImVector_DockNodeSettings
	WantFullRebuild bool
}



pub type ViewportP = C.ImGuiViewportP
@[typedef]
struct C.ImGuiViewportP {
pub mut:
	_ImGuiViewport          Viewport
	Window                  /*&Window*/voidptr= unsafe{ nil }
	Idx                     int
	LastFrameActive         int
	LastFocusedStampCount   int
	LastNameHash            ID
	LastPos                 ImVec2
	LastSize                ImVec2
	Alpha                   f32
	LastAlpha               f32
	LastFocusedHadNavWindow bool
	PlatformMonitor         i16
	BgFgDrawListsLastFrame  [2]int
	BgFgDrawLists           [2]&ImDrawList
	DrawDataP               ImDrawData
	DrawDataBuilder         ImDrawDataBuilder
	LastPlatformPos         ImVec2
	LastPlatformSize        ImVec2
	LastRendererSize        ImVec2
	WorkInsetMin            ImVec2
	WorkInsetMax            ImVec2
	BuildWorkInsetMin       ImVec2
	BuildWorkInsetMax       ImVec2
}



pub type WindowSettings = C.ImGuiWindowSettings
@[typedef]
struct C.ImGuiWindowSettings {
pub mut:
	ID          ID
	Pos         ImVec2ih
	Size        ImVec2ih
	ViewportPos ImVec2ih
	ViewportId  ID
	DockId      ID
	ClassId     ID
	DockOrder   i16
	Collapsed   bool
	IsChild     bool
	WantApply   bool
	WantDelete  bool
}



pub type SettingsHandler = C.ImGuiSettingsHandler
@[typedef]
struct C.ImGuiSettingsHandler {
pub mut:
	TypeName   /*&i8*/voidptr= unsafe{ nil }
	TypeHash   ID
	ClearAllFn fn (&Context, &SettingsHandler)
	ReadInitFn fn (&Context, &SettingsHandler)
	ReadOpenFn fn (&Context, &SettingsHandler, &i8) voidptr
	ReadLineFn fn (&Context, &SettingsHandler, voidptr, &i8)
	ApplyAllFn fn (&Context, &SettingsHandler)
	WriteAllFn fn (&Context, &SettingsHandler, &TextBuffer)
	UserData   voidptr = unsafe{ nil }
}

enum LocKey {
 version_str                         = 0
 table_size_one                      = 1
 table_size_all_fit                  = 2
 table_size_all_default              = 3
 table_reset_order                   = 4
 windowing_main_menu_bar             = 5
 windowing_popup                     = 6
 windowing_untitled                  = 7
 open_link_s                         = 8
 copy_link                           = 9
 docking_hide_tab_bar                = 10
 docking_hold_shift_to_dock          = 11
 docking_drag_to_undock_or_move_node = 12
 count                               = 13
}



pub type LocEntry = C.ImGuiLocEntry
@[typedef]
struct C.ImGuiLocEntry {
pub mut:
	Key  LocKey
	Text /*&i8*/voidptr= unsafe{ nil }
}

type ErrorCallback = fn (&Context, voidptr, &i8)

enum DebugLogFlags_ {
 none                  = 0
 event_error           = 1 << 0
 event_active_id       = 1 << 1
 event_focus           = 1 << 2
 event_popup           = 1 << 3
 event_nav             = 1 << 4
 event_clipper         = 1 << 5
 event_selection       = 1 << 6
 event_io              = 1 << 7
 event_font            = 1 << 8
 event_input_routing   = 1 << 9
 event_docking         = 1 << 10
 event_viewport        = 1 << 11
 event_mask_           = 1 << 0 | 1 << 1 | 1 << 2 | 1 << 3 | 1 << 4 | 1 << 5 | 1 << 6 | 1 << 7 | 1 << 8 | 1 << 9 | 1 << 10 | 1 << 11
 output_to_tty         = 1 << 20
 output_to_test_engine = 1 << 21
}



pub type DebugAllocEntry = C.ImGuiDebugAllocEntry
@[typedef]
struct C.ImGuiDebugAllocEntry {
pub mut:
	FrameCount int
	AllocCount ImS16
	FreeCount  ImS16
}



pub type DebugAllocInfo = C.ImGuiDebugAllocInfo
@[typedef]
struct C.ImGuiDebugAllocInfo {
pub mut:
	TotalAllocCount int
	TotalFreeCount  int
	LastEntriesIdx  ImS16
	LastEntriesBuf  [6]DebugAllocEntry
}



pub type MetricsConfig = C.ImGuiMetricsConfig
@[typedef]
struct C.ImGuiMetricsConfig {
pub mut:
	ShowDebugLog             bool
	ShowIDStackTool          bool
	ShowWindowsRects         bool
	ShowWindowsBeginOrder    bool
	ShowTablesRects          bool
	ShowDrawCmdMesh          bool
	ShowDrawCmdBoundingBoxes bool
	ShowTextEncodingViewer   bool
	ShowDockingNodes         bool
	ShowWindowsRectsType     int
	ShowTablesRectsType      int
	HighlightMonitorIdx      int
	HighlightViewportID      ID
}



pub type StackLevelInfo = C.ImGuiStackLevelInfo
@[typedef]
struct C.ImGuiStackLevelInfo {
pub mut:
	ID              ID
	QueryFrameCount ImS8
	QuerySuccess    bool
	DataType        DataType
	Desc            [57]i8
}



pub type ImVector_StackLevelInfo = C.ImVector_ImGuiStackLevelInfo
@[typedef]
struct C.ImVector_ImGuiStackLevelInfo {
pub mut:
	Size     int
	Capacity int
	Data     /*&StackLevelInfo*/voidptr= unsafe{ nil }
}



pub type IDStackTool = C.ImGuiIDStackTool
@[typedef]
struct C.ImGuiIDStackTool {
pub mut:
	LastActiveFrame         int
	StackLevel              int
	QueryId                 ID
	Results                 ImVector_StackLevelInfo
	CopyToClipboardOnCtrlC  bool
	CopyToClipboardLastTime f32
	ResultPathBuf           TextBuffer
}

type ContextHookCallback = fn (&Context, &ContextHook)

enum ContextHookType {
 new_frame_pre
 new_frame_post
 end_frame_pre
 end_frame_post
 render_pre
 render_post
 shutdown
 pending_removal_
}



pub type ContextHook = C.ImGuiContextHook
@[typedef]
struct C.ImGuiContextHook {
pub mut:
	HookId   ID
	Type     ContextHookType
	Owner    ID
	Callback /*ContextHookCallback*/voidptr = unsafe{ nil }
	UserData voidptr = unsafe{ nil }
}



pub type ImVector_InputEvent = C.ImVector_ImGuiInputEvent
@[typedef]
struct C.ImVector_ImGuiInputEvent {
pub mut:
	Size     int
	Capacity int
	Data     /*&InputEvent*/voidptr= unsafe{ nil }
}



pub type ImVector_WindowStackData = C.ImVector_ImGuiWindowStackData
@[typedef]
struct C.ImVector_ImGuiWindowStackData {
pub mut:
	Size     int
	Capacity int
	Data     /*&WindowStackData*/voidptr= unsafe{ nil }
}



pub type ImVector_ColorMod = C.ImVector_ImGuiColorMod
@[typedef]
struct C.ImVector_ImGuiColorMod {
pub mut:
	Size     int
	Capacity int
	Data     /*&ColorMod*/voidptr= unsafe{ nil }
}



pub type ImVector_StyleMod = C.ImVector_ImGuiStyleMod
@[typedef]
struct C.ImVector_ImGuiStyleMod {
pub mut:
	Size     int
	Capacity int
	Data     /*&StyleMod*/voidptr= unsafe{ nil }
}



pub type ImVector_FocusScopeData = C.ImVector_ImGuiFocusScopeData
@[typedef]
struct C.ImVector_ImGuiFocusScopeData {
pub mut:
	Size     int
	Capacity int
	Data     /*&FocusScopeData*/voidptr= unsafe{ nil }
}



pub type ImVector_ItemFlags = C.ImVector_ImGuiItemFlags
@[typedef]
struct C.ImVector_ImGuiItemFlags {
pub mut:
	Size     int
	Capacity int
	Data     /*&ItemFlags*/voidptr= unsafe{ nil }
}



pub type ImVector_GroupData = C.ImVector_ImGuiGroupData
@[typedef]
struct C.ImVector_ImGuiGroupData {
pub mut:
	Size     int
	Capacity int
	Data     /*&GroupData*/voidptr= unsafe{ nil }
}



pub type ImVector_PopupData = C.ImVector_ImGuiPopupData
@[typedef]
struct C.ImVector_ImGuiPopupData {
pub mut:
	Size     int
	Capacity int
	Data     /*&PopupData*/voidptr= unsafe{ nil }
}



pub type ImVector_TreeNodeStackData = C.ImVector_ImGuiTreeNodeStackData
@[typedef]
struct C.ImVector_ImGuiTreeNodeStackData {
pub mut:
	Size     int
	Capacity int
	Data     /*&TreeNodeStackData*/voidptr= unsafe{ nil }
}



pub type ImVector_ViewportPPtr = C.ImVector_ImGuiViewportPPtr
@[typedef]
struct C.ImVector_ImGuiViewportPPtr {
pub mut:
	Size     int
	Capacity int
	Data     /*&&ViewportP*/voidptr= unsafe{ nil }
}



pub type ImVector_unsigned_char = C.ImVector_unsigned_char
@[typedef]
struct C.ImVector_unsigned_char {
pub mut:
	Size     int
	Capacity int
	Data     /*&u8*/voidptr= unsafe{ nil }
}



pub type ImVector_ListClipperData = C.ImVector_ImGuiListClipperData
@[typedef]
struct C.ImVector_ImGuiListClipperData {
pub mut:
	Size     int
	Capacity int
	Data     /*&ListClipperData*/voidptr= unsafe{ nil }
}



pub type ImVector_TableTempData = C.ImVector_ImGuiTableTempData
@[typedef]
struct C.ImVector_ImGuiTableTempData {
pub mut:
	Size     int
	Capacity int
	Data     /*&TableTempData*/voidptr= unsafe{ nil }
}



pub type ImVector_Table = C.ImVector_ImGuiTable
@[typedef]
struct C.ImVector_ImGuiTable {
pub mut:
	Size     int
	Capacity int
	Data     /*&Table*/voidptr= unsafe{ nil }
}



pub type ImPool_Table = C.ImPool_ImGuiTable
@[typedef]
struct C.ImPool_ImGuiTable {
pub mut:
	Buf        ImVector_Table
	Map        Storage
	FreeIdx    ImPoolIdx
	AliveCount ImPoolIdx
}



pub type ImVector_TabBar = C.ImVector_ImGuiTabBar
@[typedef]
struct C.ImVector_ImGuiTabBar {
pub mut:
	Size     int
	Capacity int
	Data     /*&TabBar*/voidptr= unsafe{ nil }
}



pub type ImPool_TabBar = C.ImPool_ImGuiTabBar
@[typedef]
struct C.ImPool_ImGuiTabBar {
pub mut:
	Buf        ImVector_TabBar
	Map        Storage
	FreeIdx    ImPoolIdx
	AliveCount ImPoolIdx
}



pub type ImVector_PtrOrIndex = C.ImVector_ImGuiPtrOrIndex
@[typedef]
struct C.ImVector_ImGuiPtrOrIndex {
pub mut:
	Size     int
	Capacity int
	Data     /*&PtrOrIndex*/voidptr= unsafe{ nil }
}



pub type ImVector_ShrinkWidthItem = C.ImVector_ImGuiShrinkWidthItem
@[typedef]
struct C.ImVector_ImGuiShrinkWidthItem {
pub mut:
	Size     int
	Capacity int
	Data     /*&ShrinkWidthItem*/voidptr= unsafe{ nil }
}



pub type ImVector_MultiSelectTempData = C.ImVector_ImGuiMultiSelectTempData
@[typedef]
struct C.ImVector_ImGuiMultiSelectTempData {
pub mut:
	Size     int
	Capacity int
	Data     /*&MultiSelectTempData*/voidptr= unsafe{ nil }
}



pub type ImVector_MultiSelectState = C.ImVector_ImGuiMultiSelectState
@[typedef]
struct C.ImVector_ImGuiMultiSelectState {
pub mut:
	Size     int
	Capacity int
	Data     /*&MultiSelectState*/voidptr= unsafe{ nil }
}



pub type ImPool_MultiSelectState = C.ImPool_ImGuiMultiSelectState
@[typedef]
struct C.ImPool_ImGuiMultiSelectState {
pub mut:
	Buf        ImVector_MultiSelectState
	Map        Storage
	FreeIdx    ImPoolIdx
	AliveCount ImPoolIdx
}



pub type ImVector_ID = C.ImVector_ImGuiID
@[typedef]
struct C.ImVector_ImGuiID {
pub mut:
	Size     int
	Capacity int
	Data     /*&ID*/voidptr= unsafe{ nil }
}



pub type ImVector_SettingsHandler = C.ImVector_ImGuiSettingsHandler
@[typedef]
struct C.ImVector_ImGuiSettingsHandler {
pub mut:
	Size     int
	Capacity int
	Data     /*&SettingsHandler*/voidptr= unsafe{ nil }
}



pub type ImChunkStream_WindowSettings = C.ImChunkStream_ImGuiWindowSettings
@[typedef]
struct C.ImChunkStream_ImGuiWindowSettings {
pub mut:
	Buf ImVector_char
}



pub type ImChunkStream_TableSettings = C.ImChunkStream_ImGuiTableSettings
@[typedef]
struct C.ImChunkStream_ImGuiTableSettings {
pub mut:
	Buf ImVector_char
}



pub type ImVector_ContextHook = C.ImVector_ImGuiContextHook
@[typedef]
struct C.ImVector_ImGuiContextHook {
pub mut:
	Size     int
	Capacity int
	Data     /*&ContextHook*/voidptr= unsafe{ nil }
}



pub type Context = C.ImGuiContext
@[typedef]
struct C.ImGuiContext {
pub mut:
	Initialized                        bool
	FontAtlasOwnedByContext            bool
	IO                                 IO
	PlatformIO                         PlatformIO
	Style                              Style
	ConfigFlagsCurrFrame               ConfigFlags
	ConfigFlagsLastFrame               ConfigFlags
	Font                               /*&ImFont*/voidptr= unsafe{ nil }
	FontSize                           f32
	FontBaseSize                       f32
	FontScale                          f32
	CurrentDpiScale                    f32
	DrawListSharedData                 ImDrawListSharedData
	Time                               f64
	FrameCount                         int
	FrameCountEnded                    int
	FrameCountPlatformEnded            int
	FrameCountRendered                 int
	WithinEndChildID                   ID
	WithinFrameScope                   bool
	WithinFrameScopeWithImplicitWindow bool
	GcCompactAll                       bool
	TestEngineHookItems                bool
	TestEngine                         voidptr = unsafe{ nil }
	ContextName                        [16]i8
	InputEventsQueue                   ImVector_InputEvent
	InputEventsTrail                   ImVector_InputEvent
	InputEventsNextMouseSource         MouseSource
	InputEventsNextEventId             ImU32
	Windows                            ImVector_WindowPtr
	WindowsFocusOrder                  ImVector_WindowPtr
	WindowsTempSortBuffer              ImVector_WindowPtr
	CurrentWindowStack                 ImVector_WindowStackData
	WindowsById                        Storage
	WindowsActiveCount                 int
	WindowsBorderHoverPadding          f32
	DebugBreakInWindow                 ID
	CurrentWindow                      /*&Window*/voidptr= unsafe{ nil }
	HoveredWindow                      /*&Window*/voidptr= unsafe{ nil }
	HoveredWindowUnderMovingWindow     /*&Window*/voidptr= unsafe{ nil }
	HoveredWindowBeforeClear           /*&Window*/voidptr= unsafe{ nil }
	MovingWindow                       /*&Window*/voidptr= unsafe{ nil }
	WheelingWindow                     /*&Window*/voidptr= unsafe{ nil }
	WheelingWindowRefMousePos          ImVec2
	WheelingWindowStartFrame           int
	WheelingWindowScrolledFrame        int
	WheelingWindowReleaseTimer         f32
	WheelingWindowWheelRemainder       ImVec2
	WheelingAxisAvg                    ImVec2
	DebugDrawIdConflicts               ID
	DebugHookIdInfo                    ID
	HoveredId                          ID
	HoveredIdPreviousFrame             ID
	HoveredIdPreviousFrameItemCount    int
	HoveredIdTimer                     f32
	HoveredIdNotActiveTimer            f32
	HoveredIdAllowOverlap              bool
	HoveredIdIsDisabled                bool
	ItemUnclipByLog                    bool
	ActiveId                           ID
	ActiveIdIsAlive                    ID
	ActiveIdTimer                      f32
	ActiveIdIsJustActivated            bool
	ActiveIdAllowOverlap               bool
	ActiveIdNoClearOnFocusLoss         bool
	ActiveIdHasBeenPressedBefore       bool
	ActiveIdHasBeenEditedBefore        bool
	ActiveIdHasBeenEditedThisFrame     bool
	ActiveIdFromShortcut               bool
	ActiveIdMouseButton                int
	ActiveIdClickOffset                ImVec2
	ActiveIdWindow                     /*&Window*/voidptr= unsafe{ nil }
	ActiveIdSource                     InputSource
	ActiveIdPreviousFrame              ID
	DeactivatedItemData                DeactivatedItemData
	ActiveIdValueOnActivation          DataTypeStorage
	LastActiveId                       ID
	LastActiveIdTimer                  f32
	LastKeyModsChangeTime              f64
	LastKeyModsChangeFromNoneTime      f64
	LastKeyboardKeyPressTime           f64
	KeysMayBeCharInput                 ImBitArrayForNamedKeys
	KeysOwnerData                      [155]KeyOwnerData
	KeysRoutingTable                   KeyRoutingTable
	ActiveIdUsingNavDirMask            ImU32
	ActiveIdUsingAllKeyboardKeys       bool
	DebugBreakInShortcutRouting        KeyChord
	CurrentFocusScopeId                ID
	CurrentItemFlags                   ItemFlags
	DebugLocateId                      ID
	NextItemData                       NextItemData
	LastItemData                       LastItemData
	NextWindowData                     NextWindowData
	DebugShowGroupRects                bool
	DebugFlashStyleColorIdx            Col
	ColorStack                         ImVector_ColorMod
	StyleVarStack                      ImVector_StyleMod
	FontStack                          ImVector_ImFontPtr
	FocusScopeStack                    ImVector_FocusScopeData
	ItemFlagsStack                     ImVector_ItemFlags
	GroupStack                         ImVector_GroupData
	OpenPopupStack                     ImVector_PopupData
	BeginPopupStack                    ImVector_PopupData
	TreeNodeStack                      ImVector_TreeNodeStackData
	Viewports                          ImVector_ViewportPPtr
	CurrentViewport                    /*&ViewportP*/voidptr= unsafe{ nil }
	MouseViewport                      /*&ViewportP*/voidptr= unsafe{ nil }
	MouseLastHoveredViewport           /*&ViewportP*/voidptr= unsafe{ nil }
	PlatformLastFocusedViewportId      ID
	FallbackMonitor                    PlatformMonitor
	PlatformMonitorsFullWorkRect       ImRect
	ViewportCreatedCount               int
	PlatformWindowsCreatedCount        int
	ViewportFocusedStampCount          int
	NavCursorVisible                   bool
	NavHighlightItemUnderNav           bool
	NavMousePosDirty                   bool
	NavIdIsAlive                       bool
	NavId                              ID
	NavWindow                          /*&Window*/voidptr= unsafe{ nil }
	NavFocusScopeId                    ID
	NavLayer                           NavLayer
	NavActivateId                      ID
	NavActivateDownId                  ID
	NavActivatePressedId               ID
	NavActivateFlags                   ActivateFlags
	NavFocusRoute                      ImVector_FocusScopeData
	NavHighlightActivatedId            ID
	NavHighlightActivatedTimer         f32
	NavNextActivateId                  ID
	NavNextActivateFlags               ActivateFlags
	NavInputSource                     InputSource
	NavLastValidSelectionUserData      SelectionUserData
	NavCursorHideFrames                ImS8
	NavAnyRequest                      bool
	NavInitRequest                     bool
	NavInitRequestFromMove             bool
	NavInitResult                      NavItemData
	NavMoveSubmitted                   bool
	NavMoveScoringItems                bool
	NavMoveForwardToNextFrame          bool
	NavMoveFlags                       NavMoveFlags
	NavMoveScrollFlags                 ScrollFlags
	NavMoveKeyMods                     KeyChord
	NavMoveDir                         Dir
	NavMoveDirForDebug                 Dir
	NavMoveClipDir                     Dir
	NavScoringRect                     ImRect
	NavScoringNoClipRect               ImRect
	NavScoringDebugCount               int
	NavTabbingDir                      int
	NavTabbingCounter                  int
	NavMoveResultLocal                 NavItemData
	NavMoveResultLocalVisible          NavItemData
	NavMoveResultOther                 NavItemData
	NavTabbingResultFirst              NavItemData
	NavJustMovedFromFocusScopeId       ID
	NavJustMovedToId                   ID
	NavJustMovedToFocusScopeId         ID
	NavJustMovedToKeyMods              KeyChord
	NavJustMovedToIsTabbing            bool
	NavJustMovedToHasSelectionData     bool
	ConfigNavWindowingKeyNext          KeyChord
	ConfigNavWindowingKeyPrev          KeyChord
	NavWindowingTarget                 /*&Window*/voidptr= unsafe{ nil }
	NavWindowingTargetAnim             /*&Window*/voidptr= unsafe{ nil }
	NavWindowingListWindow             /*&Window*/voidptr= unsafe{ nil }
	NavWindowingTimer                  f32
	NavWindowingHighlightAlpha         f32
	NavWindowingToggleLayer            bool
	NavWindowingToggleKey              Key
	NavWindowingAccumDeltaPos          ImVec2
	NavWindowingAccumDeltaSize         ImVec2
	DimBgRatio                         f32
	DragDropActive                     bool
	DragDropWithinSource               bool
	DragDropWithinTarget               bool
	DragDropSourceFlags                DragDropFlags
	DragDropSourceFrameCount           int
	DragDropMouseButton                int
	DragDropPayload                    Payload
	DragDropTargetRect                 ImRect
	DragDropTargetClipRect             ImRect
	DragDropTargetId                   ID
	DragDropAcceptFlags                DragDropFlags
	DragDropAcceptIdCurrRectSurface    f32
	DragDropAcceptIdCurr               ID
	DragDropAcceptIdPrev               ID
	DragDropAcceptFrameCount           int
	DragDropHoldJustPressedId          ID
	DragDropPayloadBufHeap             ImVector_unsigned_char
	DragDropPayloadBufLocal            [16]u8
	ClipperTempDataStacked             int
	ClipperTempData                    ImVector_ListClipperData
	CurrentTable                       /*&Table*/voidptr= unsafe{ nil }
	DebugBreakInTable                  ID
	TablesTempDataStacked              int
	TablesTempData                     ImVector_TableTempData
	Tables                             ImPool_Table
	TablesLastTimeActive               ImVector_float
	DrawChannelsTempMergeBuffer        ImVector_ImDrawChannel
	CurrentTabBar                      /*&TabBar*/voidptr= unsafe{ nil }
	TabBars                            ImPool_TabBar
	CurrentTabBarStack                 ImVector_PtrOrIndex
	ShrinkWidthBuffer                  ImVector_ShrinkWidthItem
	BoxSelectState                     BoxSelectState
	CurrentMultiSelect                 /*&MultiSelectTempData*/voidptr= unsafe{ nil }
	MultiSelectTempDataStacked         int
	MultiSelectTempData                ImVector_MultiSelectTempData
	MultiSelectStorage                 ImPool_MultiSelectState
	HoverItemDelayId                   ID
	HoverItemDelayIdPreviousFrame      ID
	HoverItemDelayTimer                f32
	HoverItemDelayClearTimer           f32
	HoverItemUnlockedStationaryId      ID
	HoverWindowUnlockedStationaryId    ID
	MouseCursor                        MouseCursor
	MouseStationaryTimer               f32
	MouseLastValidPos                  ImVec2
	InputTextState                     InputTextState
	InputTextDeactivatedState          InputTextDeactivatedState
	InputTextPasswordFont              ImFont
	TempInputId                        ID
	DataTypeZeroValue                  DataTypeStorage
	BeginMenuDepth                     int
	BeginComboDepth                    int
	ColorEditOptions                   ColorEditFlags
	ColorEditCurrentID                 ID
	ColorEditSavedID                   ID
	ColorEditSavedHue                  f32
	ColorEditSavedSat                  f32
	ColorEditSavedColor                ImU32
	ColorPickerRef                     ImVec4
	ComboPreviewData                   ComboPreviewData
	WindowResizeBorderExpectedRect     ImRect
	WindowResizeRelativeMode           bool
	ScrollbarSeekMode                  i16
	ScrollbarClickDeltaToGrabCenter    f32
	SliderGrabClickOffset              f32
	SliderCurrentAccum                 f32
	SliderCurrentAccumDirty            bool
	DragCurrentAccumDirty              bool
	DragCurrentAccum                   f32
	DragSpeedDefaultRatio              f32
	DisabledAlphaBackup                f32
	DisabledStackSize                  i16
	TooltipOverrideCount               i16
	TooltipPreviousWindow              /*&Window*/voidptr= unsafe{ nil }
	ClipboardHandlerData               ImVector_char
	MenusIdSubmittedThisFrame          ImVector_ID
	TypingSelectState                  TypingSelectState
	PlatformImeData                    PlatformImeData
	PlatformImeDataPrev                PlatformImeData
	PlatformImeViewport                ID
	DockContext                        DockContext
	DockNodeWindowMenuHandler          fn (&Context, &DockNode, &TabBar)
	SettingsLoaded                     bool
	SettingsDirtyTimer                 f32
	SettingsIniData                    TextBuffer
	SettingsHandlers                   ImVector_SettingsHandler
	SettingsWindows                    ImChunkStream_WindowSettings
	SettingsTables                     ImChunkStream_TableSettings
	Hooks                              ImVector_ContextHook
	HookIdNext                         ID
	LocalizationTable                  [13]&i8
	LogEnabled                         bool
	LogFlags                           LogFlags
	LogWindow                          /*&Window*/voidptr= unsafe{ nil }
	LogFile                            /*ImFileHandle*/voidptr = unsafe{ nil }
	LogBuffer                          TextBuffer
	LogNextPrefix                      /*&i8*/voidptr= unsafe{ nil }
	LogNextSuffix                      /*&i8*/voidptr= unsafe{ nil }
	LogLinePosY                        f32
	LogLineFirstItem                   bool
	LogDepthRef                        int
	LogDepthToExpand                   int
	LogDepthToExpandDefault            int
	ErrorCallback                      /*ErrorCallback*/voidptr = unsafe{ nil }
	ErrorCallbackUserData              voidptr = unsafe{ nil }
	ErrorTooltipLockedPos              ImVec2
	ErrorFirst                         bool
	ErrorCountCurrentFrame             int
	StackSizesInNewFrame               ErrorRecoveryState
	StackSizesInBeginForCurrentWindow  /*&ErrorRecoveryState*/voidptr= unsafe{ nil }
	DebugDrawIdConflictsCount          int
	DebugLogFlags                      DebugLogFlags
	DebugLogBuf                        TextBuffer
	DebugLogIndex                      TextIndex
	DebugLogSkippedErrors              int
	DebugLogAutoDisableFlags           DebugLogFlags
	DebugLogAutoDisableFrames          ImU8
	DebugLocateFrames                  ImU8
	DebugBreakInLocateId               bool
	DebugBreakKeyChord                 KeyChord
	DebugBeginReturnValueCullDepth     ImS8
	DebugItemPickerActive              bool
	DebugItemPickerMouseButton         ImU8
	DebugItemPickerBreakId             ID
	DebugFlashStyleColorTime           f32
	DebugFlashStyleColorBackup         ImVec4
	DebugMetricsConfig                 MetricsConfig
	DebugIDStackTool                   IDStackTool
	DebugAllocInfo                     DebugAllocInfo
	DebugHoveredDockNode               /*&DockNode*/voidptr= unsafe{ nil }
	FramerateSecPerFrame               [60]f32
	FramerateSecPerFrameIdx            int
	FramerateSecPerFrameCount          int
	FramerateSecPerFrameAccum          f32
	WantCaptureMouseNextFrame          int
	WantCaptureKeyboardNextFrame       int
	WantTextInputNextFrame             int
	TempBuffer                         ImVector_char
	TempKeychordName                   [64]i8
}



pub type WindowTempData = C.ImGuiWindowTempData
@[typedef]
struct C.ImGuiWindowTempData {
pub mut:
	CursorPos                 ImVec2
	CursorPosPrevLine         ImVec2
	CursorStartPos            ImVec2
	CursorMaxPos              ImVec2
	IdealMaxPos               ImVec2
	CurrLineSize              ImVec2
	PrevLineSize              ImVec2
	CurrLineTextBaseOffset    f32
	PrevLineTextBaseOffset    f32
	IsSameLine                bool
	IsSetPos                  bool
	Indent                    ImVec1
	ColumnsOffset             ImVec1
	GroupOffset               ImVec1
	CursorStartPosLossyness   ImVec2
	NavLayerCurrent           NavLayer
	NavLayersActiveMask       i16
	NavLayersActiveMaskNext   i16
	NavIsScrollPushableX      bool
	NavHideHighlightOneFrame  bool
	NavWindowHasScrollY       bool
	MenuBarAppending          bool
	MenuBarOffset             ImVec2
	MenuColumns               MenuColumns
	TreeDepth                 int
	TreeHasStackDataDepthMask ImU32
	ChildWindows              ImVector_WindowPtr
	StateStorage              /*&Storage*/voidptr= unsafe{ nil }
	CurrentColumns            /*&OldColumns*/voidptr= unsafe{ nil }
	CurrentTableIdx           int
	LayoutType                LayoutType
	ParentLayoutType          LayoutType
	ModalDimBgColor           ImU32
	WindowItemStatusFlags     ItemStatusFlags
	ChildItemStatusFlags      ItemStatusFlags
	DockTabItemStatusFlags    ItemStatusFlags
	DockTabItemRect           ImRect
	ItemWidth                 f32
	TextWrapPos               f32
	ItemWidthStack            ImVector_float
	TextWrapPosStack          ImVector_float
}



pub type ImVector_OldColumns = C.ImVector_ImGuiOldColumns
@[typedef]
struct C.ImVector_ImGuiOldColumns {
pub mut:
	Size     int
	Capacity int
	Data     /*&OldColumns*/voidptr= unsafe{ nil }
}



pub type Window = C.ImGuiWindow
@[typedef]
struct C.ImGuiWindow {
pub mut:
	Ctx                                /*&Context*/voidptr= unsafe{ nil }
	Name                               /*&i8*/voidptr= unsafe{ nil }
	ID                                 ID
	Flags                              WindowFlags
	FlagsPreviousFrame                 WindowFlags
	ChildFlags                         ChildFlags
	WindowClass                        WindowClass
	Viewport                           /*&ViewportP*/voidptr= unsafe{ nil }
	ViewportId                         ID
	ViewportPos                        ImVec2
	ViewportAllowPlatformMonitorExtend int
	Pos                                ImVec2
	Size                               ImVec2
	SizeFull                           ImVec2
	ContentSize                        ImVec2
	ContentSizeIdeal                   ImVec2
	ContentSizeExplicit                ImVec2
	WindowPadding                      ImVec2
	WindowRounding                     f32
	WindowBorderSize                   f32
	TitleBarHeight                     f32
	MenuBarHeight                      f32
	DecoOuterSizeX1                    f32
	DecoOuterSizeY1                    f32
	DecoOuterSizeX2                    f32
	DecoOuterSizeY2                    f32
	DecoInnerSizeX1                    f32
	DecoInnerSizeY1                    f32
	NameBufLen                         int
	MoveId                             ID
	TabId                              ID
	ChildId                            ID
	PopupId                            ID
	Scroll                             ImVec2
	ScrollMax                          ImVec2
	ScrollTarget                       ImVec2
	ScrollTargetCenterRatio            ImVec2
	ScrollTargetEdgeSnapDist           ImVec2
	ScrollbarSizes                     ImVec2
	ScrollbarX                         bool
	ScrollbarY                         bool
	ScrollbarXStabilizeEnabled         bool
	ScrollbarXStabilizeToggledHistory  ImU8
	ViewportOwned                      bool
	Active                             bool
	WasActive                          bool
	WriteAccessed                      bool
	Collapsed                          bool
	WantCollapseToggle                 bool
	SkipItems                          bool
	SkipRefresh                        bool
	Appearing                          bool
	Hidden                             bool
	IsFallbackWindow                   bool
	IsExplicitChild                    bool
	HasCloseButton                     bool
	ResizeBorderHovered                i8
	ResizeBorderHeld                   i8
	BeginCount                         i16
	BeginCountPreviousFrame            i16
	BeginOrderWithinParent             i16
	BeginOrderWithinContext            i16
	FocusOrder                         i16
	AutoFitFramesX                     ImS8
	AutoFitFramesY                     ImS8
	AutoFitOnlyGrows                   bool
	AutoPosLastDirection               Dir
	HiddenFramesCanSkipItems           ImS8
	HiddenFramesCannotSkipItems        ImS8
	HiddenFramesForRenderOnly          ImS8
	DisableInputsFrames                ImS8
	SetWindowPosAllowFlags             Cond
	SetWindowSizeAllowFlags            Cond
	SetWindowCollapsedAllowFlags       Cond
	SetWindowDockAllowFlags            Cond
	SetWindowPosVal                    ImVec2
	SetWindowPosPivot                  ImVec2
	IDStack                            ImVector_ID
	DC                                 WindowTempData
	OuterRectClipped                   ImRect
	InnerRect                          ImRect
	InnerClipRect                      ImRect
	WorkRect                           ImRect
	ParentWorkRect                     ImRect
	ClipRect                           ImRect
	ContentRegionRect                  ImRect
	HitTestHoleSize                    ImVec2ih
	HitTestHoleOffset                  ImVec2ih
	LastFrameActive                    int
	LastFrameJustFocused               int
	LastTimeActive                     f32
	ItemWidthDefault                   f32
	StateStorage                       Storage
	ColumnsStorage                     ImVector_OldColumns
	FontWindowScale                    f32
	FontWindowScaleParents             f32
	FontDpiScale                       f32
	FontRefSize                        f32
	SettingsOffset                     int
	DrawList                           /*&ImDrawList*/voidptr= unsafe{ nil }
	DrawListInst                       ImDrawList
	ParentWindow                       /*&Window*/voidptr= unsafe{ nil }
	ParentWindowInBeginStack           /*&Window*/voidptr= unsafe{ nil }
	RootWindow                         /*&Window*/voidptr= unsafe{ nil }
	RootWindowPopupTree                /*&Window*/voidptr= unsafe{ nil }
	RootWindowDockTree                 /*&Window*/voidptr= unsafe{ nil }
	RootWindowForTitleBarHighlight     /*&Window*/voidptr= unsafe{ nil }
	RootWindowForNav                   /*&Window*/voidptr= unsafe{ nil }
	ParentWindowForFocusRoute          /*&Window*/voidptr= unsafe{ nil }
	NavLastChildNavWindow              /*&Window*/voidptr= unsafe{ nil }
	NavLastIds                         [2]ID
	NavRectRel                         [2]ImRect
	NavPreferredScoringPosRel          [2]ImVec2
	NavRootFocusScopeId                ID
	MemoryDrawListIdxCapacity          int
	MemoryDrawListVtxCapacity          int
	MemoryCompacted                    bool
	DockIsActive                       bool
	DockNodeIsVisible                  bool
	DockTabIsVisible                   bool
	DockTabWantClose                   bool
	DockOrder                          i16
	DockStyle                          WindowDockStyle
	DockNode                           /*&DockNode*/voidptr= unsafe{ nil }
	DockNodeAsHost                     /*&DockNode*/voidptr= unsafe{ nil }
	DockId                             ID
}

enum TabBarFlagsPrivate_ {
 dock_node     = 1 << 20
 is_focused    = 1 << 21
 save_settings = 1 << 22
}

enum TabItemFlagsPrivate_ {
 section_mask_   = 1 << 6 | 1 << 7
 no_close_button = 1 << 20
 button          = 1 << 21
 invisible       = 1 << 22
 unsorted        = 1 << 23
}



pub type TabItem = C.ImGuiTabItem
@[typedef]
struct C.ImGuiTabItem {
pub mut:
	ID                ID
	Flags             TabItemFlags
	Window            /*&Window*/voidptr= unsafe{ nil }
	LastFrameVisible  int
	LastFrameSelected int
	Offset            f32
	Width             f32
	ContentWidth      f32
	RequestedWidth    f32
	NameOffset        ImS32
	BeginOrder        ImS16
	IndexDuringLayout ImS16
	WantClose         bool
}



pub type ImVector_TabItem = C.ImVector_ImGuiTabItem
@[typedef]
struct C.ImVector_ImGuiTabItem {
pub mut:
	Size     int
	Capacity int
	Data     /*&TabItem*/voidptr= unsafe{ nil }
}



pub type TabBar = C.ImGuiTabBar
@[typedef]
struct C.ImGuiTabBar {
pub mut:
	Window                          /*&Window*/voidptr= unsafe{ nil }
	Tabs                            ImVector_TabItem
	Flags                           TabBarFlags
	ID                              ID
	SelectedTabId                   ID
	NextSelectedTabId               ID
	VisibleTabId                    ID
	CurrFrameVisible                int
	PrevFrameVisible                int
	BarRect                         ImRect
	CurrTabsContentsHeight          f32
	PrevTabsContentsHeight          f32
	WidthAllTabs                    f32
	WidthAllTabsIdeal               f32
	ScrollingAnim                   f32
	ScrollingTarget                 f32
	ScrollingTargetDistToVisibility f32
	ScrollingSpeed                  f32
	ScrollingRectMinX               f32
	ScrollingRectMaxX               f32
	SeparatorMinX                   f32
	SeparatorMaxX                   f32
	ReorderRequestTabId             ID
	ReorderRequestOffset            ImS16
	BeginCount                      ImS8
	WantLayout                      bool
	VisibleTabWasSubmitted          bool
	TabsAddedNew                    bool
	TabsActiveCount                 ImS16
	LastTabItemIdx                  ImS16
	ItemSpacingY                    f32
	FramePadding                    ImVec2
	BackupCursorPos                 ImVec2
	TabsNames                       TextBuffer
}

type TableColumnIdx = i16
type TableDrawChannelIdx = u16



pub type TableColumn = C.ImGuiTableColumn
@[typedef]
struct C.ImGuiTableColumn {
pub mut:
	Flags                    TableColumnFlags
	WidthGiven               f32
	MinX                     f32
	MaxX                     f32
	WidthRequest             f32
	WidthAuto                f32
	WidthMax                 f32
	StretchWeight            f32
	InitStretchWeightOrWidth f32
	ClipRect                 ImRect
	UserID                   ID
	WorkMinX                 f32
	WorkMaxX                 f32
	ItemWidth                f32
	ContentMaxXFrozen        f32
	ContentMaxXUnfrozen      f32
	ContentMaxXHeadersUsed   f32
	ContentMaxXHeadersIdeal  f32
	NameOffset               ImS16
	DisplayOrder             TableColumnIdx
	IndexWithinEnabledSet    TableColumnIdx
	PrevEnabledColumn        TableColumnIdx
	NextEnabledColumn        TableColumnIdx
	SortOrder                TableColumnIdx
	DrawChannelCurrent       TableDrawChannelIdx
	DrawChannelFrozen        TableDrawChannelIdx
	DrawChannelUnfrozen      TableDrawChannelIdx
	IsEnabled                bool
	IsUserEnabled            bool
	IsUserEnabledNextFrame   bool
	IsVisibleX               bool
	IsVisibleY               bool
	IsRequestOutput          bool
	IsSkipItems              bool
	IsPreserveWidthAuto      bool
	NavLayerCurrent          ImS8
	AutoFitQueue             ImU8
	CannotSkipItemsQueue     ImU8
	SortDirection            ImU8
	SortDirectionsAvailCount ImU8
	SortDirectionsAvailMask  ImU8
	SortDirectionsAvailList  ImU8
}



pub type TableCellData = C.ImGuiTableCellData
@[typedef]
struct C.ImGuiTableCellData {
pub mut:
	BgColor ImU32
	Column  TableColumnIdx
}



pub type TableHeaderData = C.ImGuiTableHeaderData
@[typedef]
struct C.ImGuiTableHeaderData {
pub mut:
	Index     TableColumnIdx
	TextColor ImU32
	BgColor0  ImU32
	BgColor1  ImU32
}



pub type TableInstanceData = C.ImGuiTableInstanceData
@[typedef]
struct C.ImGuiTableInstanceData {
pub mut:
	TableInstanceID         ID
	LastOuterHeight         f32
	LastTopHeadersRowHeight f32
	LastFrozenHeight        f32
	HoveredRowLast          int
	HoveredRowNext          int
}



pub type ImSpan_TableColumn = C.ImSpan_ImGuiTableColumn
@[typedef]
struct C.ImSpan_ImGuiTableColumn {
pub mut:
	Data    /*&TableColumn*/voidptr= unsafe{ nil }
	DataEnd /*&TableColumn*/voidptr= unsafe{ nil }
}



pub type ImSpan_TableColumnIdx = C.ImSpan_ImGuiTableColumnIdx
@[typedef]
struct C.ImSpan_ImGuiTableColumnIdx {
pub mut:
	Data    /*&TableColumnIdx*/voidptr= unsafe{ nil }
	DataEnd /*&TableColumnIdx*/voidptr= unsafe{ nil }
}



pub type ImSpan_TableCellData = C.ImSpan_ImGuiTableCellData
@[typedef]
struct C.ImSpan_ImGuiTableCellData {
pub mut:
	Data    /*&TableCellData*/voidptr= unsafe{ nil }
	DataEnd /*&TableCellData*/voidptr= unsafe{ nil }
}



pub type ImVector_TableInstanceData = C.ImVector_ImGuiTableInstanceData
@[typedef]
struct C.ImVector_ImGuiTableInstanceData {
pub mut:
	Size     int
	Capacity int
	Data     /*&TableInstanceData*/voidptr= unsafe{ nil }
}



pub type ImVector_TableColumnSortSpecs = C.ImVector_ImGuiTableColumnSortSpecs
@[typedef]
struct C.ImVector_ImGuiTableColumnSortSpecs {
pub mut:
	Size     int
	Capacity int
	Data     /*&TableColumnSortSpecs*/voidptr= unsafe{ nil }
}



pub type Table = C.ImGuiTable
@[typedef]
struct C.ImGuiTable {
pub mut:
	ID                         ID
	Flags                      TableFlags
	RawData                    voidptr = unsafe{ nil }
	TempData                   /*&TableTempData*/voidptr= unsafe{ nil }
	Columns                    ImSpan_TableColumn
	DisplayOrderToIndex        ImSpan_TableColumnIdx
	RowCellData                ImSpan_TableCellData
	EnabledMaskByDisplayOrder  /*ImBitArrayPtr*/voidptr = unsafe{ nil }
	EnabledMaskByIndex         /*ImBitArrayPtr*/voidptr = unsafe{ nil }
	VisibleMaskByIndex         /*ImBitArrayPtr*/voidptr = unsafe{ nil }
	SettingsLoadedFlags        TableFlags
	SettingsOffset             int
	LastFrameActive            int
	ColumnsCount               int
	CurrentRow                 int
	CurrentColumn              int
	InstanceCurrent            ImS16
	InstanceInteracted         ImS16
	RowPosY1                   f32
	RowPosY2                   f32
	RowMinHeight               f32
	RowCellPaddingY            f32
	RowTextBaseline            f32
	RowIndentOffsetX           f32
	RowFlags                   TableRowFlags
	LastRowFlags               TableRowFlags
	RowBgColorCounter          int
	RowBgColor                 [2]ImU32
	BorderColorStrong          ImU32
	BorderColorLight           ImU32
	BorderX1                   f32
	BorderX2                   f32
	HostIndentX                f32
	MinColumnWidth             f32
	OuterPaddingX              f32
	CellPaddingX               f32
	CellSpacingX1              f32
	CellSpacingX2              f32
	InnerWidth                 f32
	ColumnsGivenWidth          f32
	ColumnsAutoFitWidth        f32
	ColumnsStretchSumWeights   f32
	ResizedColumnNextWidth     f32
	ResizeLockMinContentsX2    f32
	RefScale                   f32
	AngledHeadersHeight        f32
	AngledHeadersSlope         f32
	OuterRect                  ImRect
	InnerRect                  ImRect
	WorkRect                   ImRect
	InnerClipRect              ImRect
	BgClipRect                 ImRect
	Bg0ClipRectForDrawCmd      ImRect
	Bg2ClipRectForDrawCmd      ImRect
	HostClipRect               ImRect
	HostBackupInnerClipRect    ImRect
	OuterWindow                /*&Window*/voidptr= unsafe{ nil }
	InnerWindow                /*&Window*/voidptr= unsafe{ nil }
	ColumnsNames               TextBuffer
	DrawSplitter               /*&ImDrawListSplitter*/voidptr= unsafe{ nil }
	InstanceDataFirst          TableInstanceData
	InstanceDataExtra          ImVector_TableInstanceData
	SortSpecsSingle            TableColumnSortSpecs
	SortSpecsMulti             ImVector_TableColumnSortSpecs
	SortSpecs                  TableSortSpecs
	SortSpecsCount             TableColumnIdx
	ColumnsEnabledCount        TableColumnIdx
	ColumnsEnabledFixedCount   TableColumnIdx
	DeclColumnsCount           TableColumnIdx
	AngledHeadersCount         TableColumnIdx
	HoveredColumnBody          TableColumnIdx
	HoveredColumnBorder        TableColumnIdx
	HighlightColumnHeader      TableColumnIdx
	AutoFitSingleColumn        TableColumnIdx
	ResizedColumn              TableColumnIdx
	LastResizedColumn          TableColumnIdx
	HeldHeaderColumn           TableColumnIdx
	ReorderColumn              TableColumnIdx
	ReorderColumnDir           TableColumnIdx
	LeftMostEnabledColumn      TableColumnIdx
	RightMostEnabledColumn     TableColumnIdx
	LeftMostStretchedColumn    TableColumnIdx
	RightMostStretchedColumn   TableColumnIdx
	ContextPopupColumn         TableColumnIdx
	FreezeRowsRequest          TableColumnIdx
	FreezeRowsCount            TableColumnIdx
	FreezeColumnsRequest       TableColumnIdx
	FreezeColumnsCount         TableColumnIdx
	RowCellDataCurrent         TableColumnIdx
	DummyDrawChannel           TableDrawChannelIdx
	Bg2DrawChannelCurrent      TableDrawChannelIdx
	Bg2DrawChannelUnfrozen     TableDrawChannelIdx
	NavLayer                   ImS8
	IsLayoutLocked             bool
	IsInsideRow                bool
	IsInitializing             bool
	IsSortSpecsDirty           bool
	IsUsingHeaders             bool
	IsContextPopupOpen         bool
	DisableDefaultContextMenu  bool
	IsSettingsRequestLoad      bool
	IsSettingsDirty            bool
	IsDefaultDisplayOrder      bool
	IsResetAllRequest          bool
	IsResetDisplayOrderRequest bool
	IsUnfrozenRows             bool
	IsDefaultSizingPolicy      bool
	IsActiveIdAliveBeforeTable bool
	IsActiveIdInTable          bool
	HasScrollbarYCurr          bool
	HasScrollbarYPrev          bool
	MemoryCompacted            bool
	HostSkipItems              bool
}



pub type ImVector_TableHeaderData = C.ImVector_ImGuiTableHeaderData
@[typedef]
struct C.ImVector_ImGuiTableHeaderData {
pub mut:
	Size     int
	Capacity int
	Data     /*&TableHeaderData*/voidptr= unsafe{ nil }
}



pub type TableTempData = C.ImGuiTableTempData
@[typedef]
struct C.ImGuiTableTempData {
pub mut:
	TableIndex                   int
	LastTimeActive               f32
	AngledHeadersExtraWidth      f32
	AngledHeadersRequests        ImVector_TableHeaderData
	UserOuterSize                ImVec2
	DrawSplitter                 ImDrawListSplitter
	HostBackupWorkRect           ImRect
	HostBackupParentWorkRect     ImRect
	HostBackupPrevLineSize       ImVec2
	HostBackupCurrLineSize       ImVec2
	HostBackupCursorMaxPos       ImVec2
	HostBackupColumnsOffset      ImVec1
	HostBackupItemWidth          f32
	HostBackupItemWidthStackSize int
}



pub type TableColumnSettings = C.ImGuiTableColumnSettings
@[typedef]
struct C.ImGuiTableColumnSettings {
pub mut:
	WidthOrWeight f32
	UserID        ID
	Index         TableColumnIdx
	DisplayOrder  TableColumnIdx
	SortOrder     TableColumnIdx
	SortDirection ImU8
	IsEnabled     ImS8
	IsStretch     ImU8
}



pub type TableSettings = C.ImGuiTableSettings
@[typedef]
struct C.ImGuiTableSettings {
pub mut:
	ID              ID
	SaveFlags       TableFlags
	RefScale        f32
	ColumnsCount    TableColumnIdx
	ColumnsCountMax TableColumnIdx
	WantApply       bool
}



pub type ImFontBuilderIO = C.ImFontBuilderIO
@[typedef]
struct C.ImFontBuilderIO {
pub mut:
	FontBuilder_Build fn (&ImFontAtlas) bool
}

// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
// CIMGUI_DEFINE_ENUMS_AND_STRUCTS
@[c: 'ImVec2_ImVec2_Nil']
pub fn im_vec2_im_vec2_nil() &ImVec2

@[c: 'ImVec2_destroy']
pub fn im_vec2_destroy(self &ImVec2)

@[c: 'ImVec2_ImVec2_Float']
pub fn im_vec2_im_vec2_float(_x f32, _y f32) &ImVec2

@[c: 'ImVec4_ImVec4_Nil']
pub fn im_vec4_im_vec4_nil() &ImVec4

@[c: 'ImVec4_destroy']
pub fn im_vec4_destroy(self &ImVec4)

@[c: 'ImVec4_ImVec4_Float']
pub fn im_vec4_im_vec4_float(_x f32, _y f32, _z f32, _w f32) &ImVec4

@[c: 'igCreateContext']
pub fn create_context(shared_font_atlas &ImFontAtlas) &Context

@[c: 'igDestroyContext']
pub fn destroy_context(ctx &Context)

@[c: 'igGetCurrentContext']
pub fn get_current_context() &Context

@[c: 'igSetCurrentContext']
pub fn set_current_context(ctx &Context)

@[c: 'igGetIO_Nil']
pub fn get_io_nil() &IO

@[c: 'igGetPlatformIO_Nil']
pub fn get_platform_io_nil() &PlatformIO

@[c: 'igGetStyle']
pub fn get_style() &Style

@[c: 'igNewFrame']
pub fn new_frame()

@[c: 'igEndFrame']
pub fn end_frame()

@[c: 'igRender']
pub fn render()

@[c: 'igGetDrawData']
pub fn get_draw_data() &ImDrawData

@[c: 'igShowDemoWindow']
pub fn show_demo_window(p_open &bool)

@[c: 'igShowMetricsWindow']
pub fn show_metrics_window(p_open &bool)

@[c: 'igShowDebugLogWindow']
pub fn show_debug_log_window(p_open &bool)

@[c: 'igShowIDStackToolWindow']
pub fn show_ids_tack_tool_window(p_open &bool)

@[c: 'igShowAboutWindow']
pub fn show_about_window(p_open &bool)

@[c: 'igShowStyleEditor']
pub fn show_style_editor(ref &Style)

@[c: 'igShowStyleSelector']
pub fn show_style_selector(label &i8) bool

@[c: 'igShowFontSelector']
pub fn show_font_selector(label &i8)

@[c: 'igShowUserGuide']
pub fn show_user_guide()

@[c: 'igGetVersion']
pub fn get_version() &i8

@[c: 'igStyleColorsDark']
pub fn style_colors_dark(dst &Style)

@[c: 'igStyleColorsLight']
pub fn style_colors_light(dst &Style)

@[c: 'igStyleColorsClassic']
pub fn style_colors_classic(dst &Style)

@[c: 'igBegin']
pub fn begin(name &i8, p_open &bool, flags WindowFlags) bool

@[c: 'igEnd']
pub fn end()

@[c: 'igBeginChild_Str']
pub fn begin_child_str(str_id &i8, size ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c: 'igBeginChild_ID']
pub fn begin_child_id(id ID, size ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c: 'igEndChild']
pub fn end_child()

@[c: 'igIsWindowAppearing']
pub fn is_window_appearing() bool

@[c: 'igIsWindowCollapsed']
pub fn is_window_collapsed() bool

@[c: 'igIsWindowFocused']
pub fn is_window_focused(flags FocusedFlags) bool

@[c: 'igIsWindowHovered']
pub fn is_window_hovered(flags HoveredFlags) bool

@[c: 'igGetWindowDrawList']
pub fn get_window_draw_list() &ImDrawList

@[c: 'igGetWindowDpiScale']
pub fn get_window_dpi_scale() f32

@[c: 'igGetWindowPos']
pub fn get_window_pos(p_out &ImVec2)

@[c: 'igGetWindowSize']
pub fn get_window_size(p_out &ImVec2)

@[c: 'igGetWindowWidth']
pub fn get_window_width() f32

@[c: 'igGetWindowHeight']
pub fn get_window_height() f32

@[c: 'igGetWindowViewport']
pub fn get_window_viewport() &Viewport

@[c: 'igSetNextWindowPos']
pub fn set_next_window_pos(pos ImVec2, cond Cond, pivot ImVec2)

@[c: 'igSetNextWindowSize']
pub fn set_next_window_size(size ImVec2, cond Cond)

@[c: 'igSetNextWindowSizeConstraints']
pub fn set_next_window_size_constraints(size_min ImVec2, size_max ImVec2, custom_callback SizeCallback, custom_callback_data voidptr)

@[c: 'igSetNextWindowContentSize']
pub fn set_next_window_content_size(size ImVec2)

@[c: 'igSetNextWindowCollapsed']
pub fn set_next_window_collapsed(collapsed bool, cond Cond)

@[c: 'igSetNextWindowFocus']
pub fn set_next_window_focus()

@[c: 'igSetNextWindowScroll']
pub fn set_next_window_scroll(scroll ImVec2)

@[c: 'igSetNextWindowBgAlpha']
pub fn set_next_window_bg_alpha(alpha f32)

@[c: 'igSetNextWindowViewport']
pub fn set_next_window_viewport(viewport_id ID)

@[c: 'igSetWindowPos_Vec2']
pub fn set_window_pos_vec2(pos ImVec2, cond Cond)

@[c: 'igSetWindowSize_Vec2']
pub fn set_window_size_vec2(size ImVec2, cond Cond)

@[c: 'igSetWindowCollapsed_Bool']
pub fn set_window_collapsed_bool(collapsed bool, cond Cond)

@[c: 'igSetWindowFocus_Nil']
pub fn set_window_focus_nil()

@[c: 'igSetWindowFontScale']
pub fn set_window_font_scale(scale f32)

@[c: 'igSetWindowPos_Str']
pub fn set_window_pos_str(name &i8, pos ImVec2, cond Cond)

@[c: 'igSetWindowSize_Str']
pub fn set_window_size_str(name &i8, size ImVec2, cond Cond)

@[c: 'igSetWindowCollapsed_Str']
pub fn set_window_collapsed_str(name &i8, collapsed bool, cond Cond)

@[c: 'igSetWindowFocus_Str']
pub fn set_window_focus_str(name &i8)

@[c: 'igGetScrollX']
pub fn get_scroll_x() f32

@[c: 'igGetScrollY']
pub fn get_scroll_y() f32

@[c: 'igSetScrollX_Float']
pub fn set_scroll_x_float(scroll_x f32)

@[c: 'igSetScrollY_Float']
pub fn set_scroll_y_float(scroll_y f32)

@[c: 'igGetScrollMaxX']
pub fn get_scroll_max_x() f32

@[c: 'igGetScrollMaxY']
pub fn get_scroll_max_y() f32

@[c: 'igSetScrollHereX']
pub fn set_scroll_here_x(center_x_ratio f32)

@[c: 'igSetScrollHereY']
pub fn set_scroll_here_y(center_y_ratio f32)

@[c: 'igSetScrollFromPosX_Float']
pub fn set_scroll_from_pos_x_float(local_x f32, center_x_ratio f32)

@[c: 'igSetScrollFromPosY_Float']
pub fn set_scroll_from_pos_y_float(local_y f32, center_y_ratio f32)

@[c: 'igPushFont']
pub fn push_font(font &ImFont)

@[c: 'igPopFont']
pub fn pop_font()

@[c: 'igPushStyleColor_U32']
pub fn push_style_color_u32(idx Col, col ImU32)

@[c: 'igPushStyleColor_Vec4']
pub fn push_style_color_vec4(idx Col, col ImVec4)

@[c: 'igPopStyleColor']
pub fn pop_style_color(count int)

@[c: 'igPushStyleVar_Float']
pub fn push_style_var_float(idx StyleVar, val f32)

@[c: 'igPushStyleVar_Vec2']
pub fn push_style_var_vec2(idx StyleVar, val ImVec2)

@[c: 'igPushStyleVarX']
pub fn push_style_var_x(idx StyleVar, val_x f32)

@[c: 'igPushStyleVarY']
pub fn push_style_var_y(idx StyleVar, val_y f32)

@[c: 'igPopStyleVar']
pub fn pop_style_var(count int)

@[c: 'igPushItemFlag']
pub fn push_item_flag(option ItemFlags, enabled bool)

@[c: 'igPopItemFlag']
pub fn pop_item_flag()

@[c: 'igPushItemWidth']
pub fn push_item_width(item_width f32)

@[c: 'igPopItemWidth']
pub fn pop_item_width()

@[c: 'igSetNextItemWidth']
pub fn set_next_item_width(item_width f32)

@[c: 'igCalcItemWidth']
pub fn calc_item_width() f32

@[c: 'igPushTextWrapPos']
pub fn push_text_wrap_pos(wrap_local_pos_x f32)

@[c: 'igPopTextWrapPos']
pub fn pop_text_wrap_pos()

@[c: 'igGetFont']
pub fn get_font() &ImFont

@[c: 'igGetFontSize']
pub fn get_font_size() f32

@[c: 'igGetFontTexUvWhitePixel']
pub fn get_font_tex_uv_white_pixel(p_out &ImVec2)

@[c: 'igGetColorU32_Col']
pub fn get_color_u32_col(idx Col, alpha_mul f32) ImU32

@[c: 'igGetColorU32_Vec4']
pub fn get_color_u32_vec4(col ImVec4) ImU32

@[c: 'igGetColorU32_U32']
pub fn get_color_u32_u32(col ImU32, alpha_mul f32) ImU32

@[c: 'igGetStyleColorVec4']
pub fn get_style_color_vec4(idx Col) &ImVec4

@[c: 'igGetCursorScreenPos']
pub fn get_cursor_screen_pos(p_out &ImVec2)

@[c: 'igSetCursorScreenPos']
pub fn set_cursor_screen_pos(pos ImVec2)

@[c: 'igGetContentRegionAvail']
pub fn get_content_region_avail(p_out &ImVec2)

@[c: 'igGetCursorPos']
pub fn get_cursor_pos(p_out &ImVec2)

@[c: 'igGetCursorPosX']
pub fn get_cursor_pos_x() f32

@[c: 'igGetCursorPosY']
pub fn get_cursor_pos_y() f32

@[c: 'igSetCursorPos']
pub fn set_cursor_pos(local_pos ImVec2)

@[c: 'igSetCursorPosX']
pub fn set_cursor_pos_x(local_x f32)

@[c: 'igSetCursorPosY']
pub fn set_cursor_pos_y(local_y f32)

@[c: 'igGetCursorStartPos']
pub fn get_cursor_start_pos(p_out &ImVec2)

@[c: 'igSeparator']
pub fn separator()

@[c: 'igSameLine']
pub fn same_line(offset_from_start_x f32, spacing f32)

@[c: 'igNewLine']
pub fn new_line()

@[c: 'igSpacing']
pub fn spacing()

@[c: 'igDummy']
pub fn dummy(size ImVec2)

@[c: 'igIndent']
pub fn indent(indent_w f32)

@[c: 'igUnindent']
pub fn unindent(indent_w f32)

@[c: 'igBeginGroup']
pub fn begin_group()

@[c: 'igEndGroup']
pub fn end_group()

@[c: 'igAlignTextToFramePadding']
pub fn align_text_to_frame_padding()

@[c: 'igGetTextLineHeight']
pub fn get_text_line_height() f32

@[c: 'igGetTextLineHeightWithSpacing']
pub fn get_text_line_height_with_spacing() f32

@[c: 'igGetFrameHeight']
pub fn get_frame_height() f32

@[c: 'igGetFrameHeightWithSpacing']
pub fn get_frame_height_with_spacing() f32

@[c: 'igPushID_Str']
pub fn push_id_str(str_id &i8)

@[c: 'igPushID_StrStr']
pub fn push_id_str_str(str_id_begin &i8, str_id_end &i8)

@[c: 'igPushID_Ptr']
pub fn push_id_ptr(ptr_id voidptr)

@[c: 'igPushID_Int']
pub fn push_id_int(int_id int)

@[c: 'igPopID']
pub fn pop_id()

@[c: 'igGetID_Str']
pub fn get_id_str(str_id &i8) ID

@[c: 'igGetID_StrStr']
pub fn get_id_str_str(str_id_begin &i8, str_id_end &i8) ID

@[c: 'igGetID_Ptr']
pub fn get_id_ptr(ptr_id voidptr) ID

@[c: 'igGetID_Int']
pub fn get_id_int(int_id int) ID

@[c: 'igTextUnformatted']
pub fn text_unformatted(text &i8, text_end &i8)

@[c: 'igText']
@[c2v_variadic]
pub fn text(fmt ...&i8)

@[c: 'igTextV']
pub fn text_v(fmt &i8, args Va_list)

@[c: 'igTextColored']
@[c2v_variadic]
pub fn text_colored(col ImVec4, fmt ...&i8)

@[c: 'igTextColoredV']
pub fn text_colored_v(col ImVec4, fmt &i8, args Va_list)

@[c: 'igTextDisabled']
@[c2v_variadic]
pub fn text_disabled(fmt ...&i8)

@[c: 'igTextDisabledV']
pub fn text_disabled_v(fmt &i8, args Va_list)

@[c: 'igTextWrapped']
@[c2v_variadic]
pub fn text_wrapped(fmt ...&i8)

@[c: 'igTextWrappedV']
pub fn text_wrapped_v(fmt &i8, args Va_list)

@[c: 'igLabelText']
@[c2v_variadic]
pub fn label_text(label &i8, fmt ...&i8)

@[c: 'igLabelTextV']
pub fn label_text_v(label &i8, fmt &i8, args Va_list)

@[c: 'igBulletText']
@[c2v_variadic]
pub fn bullet_text(fmt ...&i8)

@[c: 'igBulletTextV']
pub fn bullet_text_v(fmt &i8, args Va_list)

@[c: 'igSeparatorText']
pub fn separator_text(label &i8)

@[c: 'igButton']
pub fn button(label &i8, size ImVec2) bool

@[c: 'igSmallButton']
pub fn small_button(label &i8) bool

@[c: 'igInvisibleButton']
pub fn invisible_button(str_id &i8, size ImVec2, flags ButtonFlags) bool

@[c: 'igArrowButton']
pub fn arrow_button(str_id &i8, dir Dir) bool

@[c: 'igCheckbox']
pub fn checkbox(label &i8, v &bool) bool

@[c: 'igCheckboxFlags_IntPtr']
pub fn checkbox_flags_int_ptr(label &i8, flags &int, flags_value int) bool

@[c: 'igCheckboxFlags_UintPtr']
pub fn checkbox_flags_uint_ptr(label &i8, flags &u32, flags_value u32) bool

@[c: 'igRadioButton_Bool']
pub fn radio_button_bool(label &i8, active bool) bool

@[c: 'igRadioButton_IntPtr']
pub fn radio_button_int_ptr(label &i8, v &int, v_button int) bool

@[c: 'igProgressBar']
pub fn progress_bar(fraction f32, size_arg ImVec2, overlay &i8)

@[c: 'igBullet']
pub fn bullet()

@[c: 'igTextLink']
pub fn text_link(label &i8) bool

@[c: 'igTextLinkOpenURL']
pub fn text_link_open_url(label &i8, url &i8)

@[c: 'igImage']
pub fn image(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2)

@[c: 'igImageWithBg']
pub fn image_with_bg(user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col ImVec4, tint_col ImVec4)

@[c: 'igImageButton']
pub fn image_button(str_id &i8, user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col ImVec4, tint_col ImVec4) bool

@[c: 'igBeginCombo']
pub fn begin_combo(label &i8, preview_value &i8, flags ComboFlags) bool

@[c: 'igEndCombo']
pub fn end_combo()

@[c: 'igCombo_Str_arr']
pub fn combo_str_arr(label &i8, current_item &int, items &&u8, items_count int, popup_max_height_in_items int) bool

@[c: 'igCombo_Str']
pub fn combo_str(label &i8, current_item &int, items_separated_by_zeros &i8, popup_max_height_in_items int) bool

@[c: 'igCombo_FnStrPtr']
pub fn combo_fn_str_ptr(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int, popup_max_height_in_items int) bool

@[c: 'igDragFloat']
pub fn drag_float(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloat2']
pub fn drag_float2(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloat3']
pub fn drag_float3(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloat4']
pub fn drag_float4(label &i8, v &f32, v_speed f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igDragFloatRange2']
pub fn drag_float_range2(label &i8, v_current_min &f32, v_current_max &f32, v_speed f32, v_min f32, v_max f32, format &i8, format_max &i8, flags SliderFlags) bool

@[c: 'igDragInt']
pub fn drag_int(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragInt2']
pub fn drag_int2(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragInt3']
pub fn drag_int3(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragInt4']
pub fn drag_int4(label &i8, v &int, v_speed f32, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igDragIntRange2']
pub fn drag_int_range2(label &i8, v_current_min &int, v_current_max &int, v_speed f32, v_min int, v_max int, format &i8, format_max &i8, flags SliderFlags) bool

@[c: 'igDragScalar']
pub fn drag_scalar(label &i8, data_type DataType, p_data voidptr, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igDragScalarN']
pub fn drag_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat']
pub fn slider_float(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat2']
pub fn slider_float2(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat3']
pub fn slider_float3(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderFloat4']
pub fn slider_float4(label &i8, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderAngle']
pub fn slider_angle(label &i8, v_rad &f32, v_degrees_min f32, v_degrees_max f32, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt']
pub fn slider_int(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt2']
pub fn slider_int2(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt3']
pub fn slider_int3(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderInt4']
pub fn slider_int4(label &i8, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igSliderScalar']
pub fn slider_scalar(label &i8, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igSliderScalarN']
pub fn slider_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igVSliderFloat']
pub fn vs_lider_float(label &i8, size ImVec2, v &f32, v_min f32, v_max f32, format &i8, flags SliderFlags) bool

@[c: 'igVSliderInt']
pub fn vs_lider_int(label &i8, size ImVec2, v &int, v_min int, v_max int, format &i8, flags SliderFlags) bool

@[c: 'igVSliderScalar']
pub fn vs_lider_scalar(label &i8, size ImVec2, data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igInputText']
pub fn input_text(label &i8, buf &i8, buf_size usize, flags InputTextFlags, callback InputTextCallback, user_data voidptr) bool

@[c: 'igInputTextMultiline']
pub fn input_text_multiline(label &i8, buf &i8, buf_size usize, size ImVec2, flags InputTextFlags, callback InputTextCallback, user_data voidptr) bool

@[c: 'igInputTextWithHint']
pub fn input_text_with_hint(label &i8, hint &i8, buf &i8, buf_size usize, flags InputTextFlags, callback InputTextCallback, user_data voidptr) bool

@[c: 'igInputFloat']
pub fn input_float(label &i8, v &f32, step f32, step_fast f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputFloat2']
pub fn input_float2(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputFloat3']
pub fn input_float3(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputFloat4']
pub fn input_float4(label &i8, v &f32, format &i8, flags InputTextFlags) bool

@[c: 'igInputInt']
pub fn input_int(label &i8, v &int, step int, step_fast int, flags InputTextFlags) bool

@[c: 'igInputInt2']
pub fn input_int2(label &i8, v &int, flags InputTextFlags) bool

@[c: 'igInputInt3']
pub fn input_int3(label &i8, v &int, flags InputTextFlags) bool

@[c: 'igInputInt4']
pub fn input_int4(label &i8, v &int, flags InputTextFlags) bool

@[c: 'igInputDouble']
pub fn input_double(label &i8, v &f64, step f64, step_fast f64, format &i8, flags InputTextFlags) bool

@[c: 'igInputScalar']
pub fn input_scalar(label &i8, data_type DataType, p_data voidptr, p_step voidptr, p_step_fast voidptr, format &i8, flags InputTextFlags) bool

@[c: 'igInputScalarN']
pub fn input_scalar_n(label &i8, data_type DataType, p_data voidptr, components int, p_step voidptr, p_step_fast voidptr, format &i8, flags InputTextFlags) bool

@[c: 'igColorEdit3']
pub fn color_edit3(label &i8, col &f32, flags ColorEditFlags) bool

@[c: 'igColorEdit4']
pub fn color_edit4(label &i8, col &f32, flags ColorEditFlags) bool

@[c: 'igColorPicker3']
pub fn color_picker3(label &i8, col &f32, flags ColorEditFlags) bool

@[c: 'igColorPicker4']
pub fn color_picker4(label &i8, col &f32, flags ColorEditFlags, ref_col &f32) bool

@[c: 'igColorButton']
pub fn color_button(desc_id &i8, col ImVec4, flags ColorEditFlags, size ImVec2) bool

@[c: 'igSetColorEditOptions']
pub fn set_color_edit_options(flags ColorEditFlags)

@[c: 'igTreeNode_Str']
pub fn tree_node_str(label &i8) bool

@[c: 'igTreeNode_StrStr']
@[c2v_variadic]
pub fn tree_node_str_str(str_id &i8, fmt ...&i8) bool

@[c: 'igTreeNode_Ptr']
@[c2v_variadic]
pub fn tree_node_ptr(ptr_id voidptr, fmt ...&i8) bool

@[c: 'igTreeNodeV_Str']
pub fn tree_node_v_str(str_id &i8, fmt &i8, args Va_list) bool

@[c: 'igTreeNodeV_Ptr']
pub fn tree_node_v_ptr(ptr_id voidptr, fmt &i8, args Va_list) bool

@[c: 'igTreeNodeEx_Str']
pub fn tree_node_ex_str(label &i8, flags TreeNodeFlags) bool

@[c: 'igTreeNodeEx_StrStr']
@[c2v_variadic]
pub fn tree_node_ex_str_str(str_id &i8, flags TreeNodeFlags, fmt ...&i8) bool

@[c: 'igTreeNodeEx_Ptr']
@[c2v_variadic]
pub fn tree_node_ex_ptr(ptr_id voidptr, flags TreeNodeFlags, fmt ...&i8) bool

@[c: 'igTreeNodeExV_Str']
pub fn tree_node_ex_v_str(str_id &i8, flags TreeNodeFlags, fmt &i8, args Va_list) bool

@[c: 'igTreeNodeExV_Ptr']
pub fn tree_node_ex_v_ptr(ptr_id voidptr, flags TreeNodeFlags, fmt &i8, args Va_list) bool

@[c: 'igTreePush_Str']
pub fn tree_push_str(str_id &i8)

@[c: 'igTreePush_Ptr']
pub fn tree_push_ptr(ptr_id voidptr)

@[c: 'igTreePop']
pub fn tree_pop()

@[c: 'igGetTreeNodeToLabelSpacing']
pub fn get_tree_node_to_label_spacing() f32

@[c: 'igCollapsingHeader_TreeNodeFlags']
pub fn collapsing_header_tree_node_flags(label &i8, flags TreeNodeFlags) bool

@[c: 'igCollapsingHeader_BoolPtr']
pub fn collapsing_header_bool_ptr(label &i8, p_visible &bool, flags TreeNodeFlags) bool

@[c: 'igSetNextItemOpen']
pub fn set_next_item_open(is_open bool, cond Cond)

@[c: 'igSetNextItemStorageID']
pub fn set_next_item_storage_id(storage_id ID)

@[c: 'igSelectable_Bool']
pub fn selectable_bool(label &i8, selected bool, flags SelectableFlags, size ImVec2) bool

@[c: 'igSelectable_BoolPtr']
pub fn selectable_bool_ptr(label &i8, p_selected &bool, flags SelectableFlags, size ImVec2) bool

@[c: 'igBeginMultiSelect']
pub fn begin_multi_select(flags MultiSelectFlags, selection_size int, items_count int) &MultiSelectIO

@[c: 'igEndMultiSelect']
pub fn end_multi_select() &MultiSelectIO

@[c: 'igSetNextItemSelectionUserData']
pub fn set_next_item_selection_user_data(selection_user_data SelectionUserData)

@[c: 'igIsItemToggledSelection']
pub fn is_item_toggled_selection() bool

@[c: 'igBeginListBox']
pub fn begin_list_box(label &i8, size ImVec2) bool

@[c: 'igEndListBox']
pub fn end_list_box()

@[c: 'igListBox_Str_arr']
pub fn list_box_str_arr(label &i8, current_item &int, items &&u8, items_count int, height_in_items int) bool

@[c: 'igListBox_FnStrPtr']
pub fn list_box_fn_str_ptr(label &i8, current_item &int, getter fn (voidptr, int) &i8, user_data voidptr, items_count int, height_in_items int) bool

@[c: 'igPlotLines_FloatPtr']
pub fn plot_lines_float_ptr(label &i8, values &f32, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2, stride int)

@[c: 'igPlotLines_FnFloatPtr']
pub fn plot_lines_fn_float_ptr(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2)

@[c: 'igPlotHistogram_FloatPtr']
pub fn plot_histogram_float_ptr(label &i8, values &f32, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2, stride int)

@[c: 'igPlotHistogram_FnFloatPtr']
pub fn plot_histogram_fn_float_ptr(label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, graph_size ImVec2)

@[c: 'igValue_Bool']
pub fn value_bool(prefix &i8, b bool)

@[c: 'igValue_Int']
pub fn value_int(prefix &i8, v int)

@[c: 'igValue_Uint']
pub fn value_uint(prefix &i8, v u32)

@[c: 'igValue_Float']
pub fn value_float(prefix &i8, v f32, float_format &i8)

@[c: 'igBeginMenuBar']
pub fn begin_menu_bar() bool

@[c: 'igEndMenuBar']
pub fn end_menu_bar()

@[c: 'igBeginMainMenuBar']
pub fn begin_main_menu_bar() bool

@[c: 'igEndMainMenuBar']
pub fn end_main_menu_bar()

@[c: 'igBeginMenu']
pub fn begin_menu(label &i8, enabled bool) bool

@[c: 'igEndMenu']
pub fn end_menu()

@[c: 'igMenuItem_Bool']
pub fn menu_item_bool(label &i8, shortcut &i8, selected bool, enabled bool) bool

@[c: 'igMenuItem_BoolPtr']
pub fn menu_item_bool_ptr(label &i8, shortcut &i8, p_selected &bool, enabled bool) bool

@[c: 'igBeginTooltip']
pub fn begin_tooltip() bool

@[c: 'igEndTooltip']
pub fn end_tooltip()

@[c: 'igSetTooltip']
@[c2v_variadic]
pub fn set_tooltip(fmt ...&i8)

@[c: 'igSetTooltipV']
pub fn set_tooltip_v(fmt &i8, args Va_list)

@[c: 'igBeginItemTooltip']
pub fn begin_item_tooltip() bool

@[c: 'igSetItemTooltip']
@[c2v_variadic]
pub fn set_item_tooltip(fmt ...&i8)

@[c: 'igSetItemTooltipV']
pub fn set_item_tooltip_v(fmt &i8, args Va_list)

@[c: 'igBeginPopup']
pub fn begin_popup(str_id &i8, flags WindowFlags) bool

@[c: 'igBeginPopupModal']
pub fn begin_popup_modal(name &i8, p_open &bool, flags WindowFlags) bool

@[c: 'igEndPopup']
pub fn end_popup()

@[c: 'igOpenPopup_Str']
pub fn open_popup_str(str_id &i8, popup_flags PopupFlags)

@[c: 'igOpenPopup_ID']
pub fn open_popup_id(id ID, popup_flags PopupFlags)

@[c: 'igOpenPopupOnItemClick']
pub fn open_popup_on_item_click(str_id &i8, popup_flags PopupFlags)

@[c: 'igCloseCurrentPopup']
pub fn close_current_popup()

@[c: 'igBeginPopupContextItem']
pub fn begin_popup_context_item(str_id &i8, popup_flags PopupFlags) bool

@[c: 'igBeginPopupContextWindow']
pub fn begin_popup_context_window(str_id &i8, popup_flags PopupFlags) bool

@[c: 'igBeginPopupContextVoid']
pub fn begin_popup_context_void(str_id &i8, popup_flags PopupFlags) bool

@[c: 'igIsPopupOpen_Str']
pub fn is_popup_open_str(str_id &i8, flags PopupFlags) bool

@[c: 'igBeginTable']
pub fn begin_table(str_id &i8, columns int, flags TableFlags, outer_size ImVec2, inner_width f32) bool

@[c: 'igEndTable']
pub fn end_table()

@[c: 'igTableNextRow']
pub fn table_next_row(row_flags TableRowFlags, min_row_height f32)

@[c: 'igTableNextColumn']
pub fn table_next_column() bool

@[c: 'igTableSetColumnIndex']
pub fn table_set_column_index(column_n int) bool

@[c: 'igTableSetupColumn']
pub fn table_setup_column(label &i8, flags TableColumnFlags, init_width_or_weight f32, user_id ID)

@[c: 'igTableSetupScrollFreeze']
pub fn table_setup_scroll_freeze(cols int, rows int)

@[c: 'igTableHeader']
pub fn table_header(label &i8)

@[c: 'igTableHeadersRow']
pub fn table_headers_row()

@[c: 'igTableAngledHeadersRow']
pub fn table_angled_headers_row()

@[c: 'igTableGetSortSpecs']
pub fn table_get_sort_specs() &TableSortSpecs

@[c: 'igTableGetColumnCount']
pub fn table_get_column_count() int

@[c: 'igTableGetColumnIndex']
pub fn table_get_column_index() int

@[c: 'igTableGetRowIndex']
pub fn table_get_row_index() int

@[c: 'igTableGetColumnName_Int']
pub fn table_get_column_name_int(column_n int) &i8

@[c: 'igTableGetColumnFlags']
pub fn table_get_column_flags(column_n int) TableColumnFlags

@[c: 'igTableSetColumnEnabled']
pub fn table_set_column_enabled(column_n int, v bool)

@[c: 'igTableGetHoveredColumn']
pub fn table_get_hovered_column() int

@[c: 'igTableSetBgColor']
pub fn table_set_bg_color(target TableBgTarget, color ImU32, column_n int)

@[c: 'igColumns']
pub fn columns(count int, id &i8, borders bool)

@[c: 'igNextColumn']
pub fn next_column()

@[c: 'igGetColumnIndex']
pub fn get_column_index() int

@[c: 'igGetColumnWidth']
pub fn get_column_width(column_index int) f32

@[c: 'igSetColumnWidth']
pub fn set_column_width(column_index int, width f32)

@[c: 'igGetColumnOffset']
pub fn get_column_offset(column_index int) f32

@[c: 'igSetColumnOffset']
pub fn set_column_offset(column_index int, offset_x f32)

@[c: 'igGetColumnsCount']
pub fn get_columns_count() int

@[c: 'igBeginTabBar']
pub fn begin_tab_bar(str_id &i8, flags TabBarFlags) bool

@[c: 'igEndTabBar']
pub fn end_tab_bar()

@[c: 'igBeginTabItem']
pub fn begin_tab_item(label &i8, p_open &bool, flags TabItemFlags) bool

@[c: 'igEndTabItem']
pub fn end_tab_item()

@[c: 'igTabItemButton']
pub fn tab_item_button(label &i8, flags TabItemFlags) bool

@[c: 'igSetTabItemClosed']
pub fn set_tab_item_closed(tab_or_docked_window_label &i8)

@[c: 'igDockSpace']
pub fn dock_space(dockspace_id ID, size ImVec2, flags DockNodeFlags, window_class &WindowClass) ID

@[c: 'igDockSpaceOverViewport']
pub fn dock_space_over_viewport(dockspace_id ID, viewport &Viewport, flags DockNodeFlags, window_class &WindowClass) ID

@[c: 'igSetNextWindowDockID']
pub fn set_next_window_dock_id(dock_id ID, cond Cond)

@[c: 'igSetNextWindowClass']
pub fn set_next_window_class(window_class &WindowClass)

@[c: 'igGetWindowDockID']
pub fn get_window_dock_id() ID

@[c: 'igIsWindowDocked']
pub fn is_window_docked() bool

@[c: 'igLogToTTY']
pub fn log_to_tty(auto_open_depth int)

@[c: 'igLogToFile']
pub fn log_to_file(auto_open_depth int, filename &i8)

@[c: 'igLogToClipboard']
pub fn log_to_clipboard(auto_open_depth int)

@[c: 'igLogFinish']
pub fn log_finish()

@[c: 'igLogButtons']
pub fn log_buttons()

@[c: 'igLogTextV']
pub fn log_text_v(fmt &i8, args Va_list)

@[c: 'igBeginDragDropSource']
pub fn begin_drag_drop_source(flags DragDropFlags) bool

@[c: 'igSetDragDropPayload']
pub fn set_drag_drop_payload(type_ &i8, data voidptr, sz usize, cond Cond) bool

@[c: 'igEndDragDropSource']
pub fn end_drag_drop_source()

@[c: 'igBeginDragDropTarget']
pub fn begin_drag_drop_target() bool

@[c: 'igAcceptDragDropPayload']
pub fn accept_drag_drop_payload(type_ &i8, flags DragDropFlags) &Payload

@[c: 'igEndDragDropTarget']
pub fn end_drag_drop_target()

@[c: 'igGetDragDropPayload']
pub fn get_drag_drop_payload() &Payload

@[c: 'igBeginDisabled']
pub fn begin_disabled(disabled bool)

@[c: 'igEndDisabled']
pub fn end_disabled()

@[c: 'igPushClipRect']
pub fn push_clip_rect(clip_rect_min ImVec2, clip_rect_max ImVec2, intersect_with_current_clip_rect bool)

@[c: 'igPopClipRect']
pub fn pop_clip_rect()

@[c: 'igSetItemDefaultFocus']
pub fn set_item_default_focus()

@[c: 'igSetKeyboardFocusHere']
pub fn set_keyboard_focus_here(offset int)

@[c: 'igSetNavCursorVisible']
pub fn set_nav_cursor_visible(visible bool)

@[c: 'igSetNextItemAllowOverlap']
pub fn set_next_item_allow_overlap()

@[c: 'igIsItemHovered']
pub fn is_item_hovered(flags HoveredFlags) bool

@[c: 'igIsItemActive']
pub fn is_item_active() bool

@[c: 'igIsItemFocused']
pub fn is_item_focused() bool

@[c: 'igIsItemClicked']
pub fn is_item_clicked(mouse_button MouseButton) bool

@[c: 'igIsItemVisible']
pub fn is_item_visible() bool

@[c: 'igIsItemEdited']
pub fn is_item_edited() bool

@[c: 'igIsItemActivated']
pub fn is_item_activated() bool

@[c: 'igIsItemDeactivated']
pub fn is_item_deactivated() bool

@[c: 'igIsItemDeactivatedAfterEdit']
pub fn is_item_deactivated_after_edit() bool

@[c: 'igIsItemToggledOpen']
pub fn is_item_toggled_open() bool

@[c: 'igIsAnyItemHovered']
pub fn is_any_item_hovered() bool

@[c: 'igIsAnyItemActive']
pub fn is_any_item_active() bool

@[c: 'igIsAnyItemFocused']
pub fn is_any_item_focused() bool

@[c: 'igGetItemID']
pub fn get_item_id() ID

@[c: 'igGetItemRectMin']
pub fn get_item_rect_min(p_out &ImVec2)

@[c: 'igGetItemRectMax']
pub fn get_item_rect_max(p_out &ImVec2)

@[c: 'igGetItemRectSize']
pub fn get_item_rect_size(p_out &ImVec2)

@[c: 'igGetMainViewport']
pub fn get_main_viewport() &Viewport

@[c: 'igGetBackgroundDrawList']
pub fn get_background_draw_list(viewport &Viewport) &ImDrawList

@[c: 'igGetForegroundDrawList_ViewportPtr']
pub fn get_foreground_draw_list_viewport_ptr(viewport &Viewport) &ImDrawList

@[c: 'igIsRectVisible_Nil']
pub fn is_rect_visible_nil(size ImVec2) bool

@[c: 'igIsRectVisible_Vec2']
pub fn is_rect_visible_vec2(rect_min ImVec2, rect_max ImVec2) bool

@[c: 'igGetTime']
pub fn get_time() f64

@[c: 'igGetFrameCount']
pub fn get_frame_count() int

@[c: 'igGetDrawListSharedData']
pub fn get_draw_list_shared_data() &ImDrawListSharedData

@[c: 'igGetStyleColorName']
pub fn get_style_color_name(idx Col) &i8

@[c: 'igSetStateStorage']
pub fn set_state_storage(storage &Storage)

@[c: 'igGetStateStorage']
pub fn get_state_storage() &Storage

@[c: 'igCalcTextSize']
pub fn calc_text_size(p_out &ImVec2, text &i8, text_end &i8, hide_text_after_double_hash bool, wrap_width f32)

@[c: 'igColorConvertU32ToFloat4']
pub fn color_convert_u32_to_float4(p_out &ImVec4, in_ ImU32)

@[c: 'igColorConvertFloat4ToU32']
pub fn color_convert_float4_to_u32(in_ ImVec4) ImU32

@[c: 'igColorConvertRGBtoHSV']
pub fn color_convert_rgb_to_hsv(r f32, g f32, b f32, out_h &f32, out_s &f32, out_v &f32)

@[c: 'igColorConvertHSVtoRGB']
pub fn color_convert_hsv_to_rgb(h f32, s f32, v f32, out_r &f32, out_g &f32, out_b &f32)

@[c: 'igIsKeyDown_Nil']
pub fn is_key_down_nil(key Key) bool

@[c: 'igIsKeyPressed_Bool']
pub fn is_key_pressed_bool(key Key, repeat bool) bool

@[c: 'igIsKeyReleased_Nil']
pub fn is_key_released_nil(key Key) bool

@[c: 'igIsKeyChordPressed_Nil']
pub fn is_key_chord_pressed_nil(key_chord KeyChord) bool

@[c: 'igGetKeyPressedAmount']
pub fn get_key_pressed_amount(key Key, repeat_delay f32, rate f32) int

@[c: 'igGetKeyName']
pub fn get_key_name(key Key) &i8

@[c: 'igSetNextFrameWantCaptureKeyboard']
pub fn set_next_frame_want_capture_keyboard(want_capture_keyboard bool)

@[c: 'igShortcut_Nil']
pub fn shortcut_nil(key_chord KeyChord, flags InputFlags) bool

@[c: 'igSetNextItemShortcut']
pub fn set_next_item_shortcut(key_chord KeyChord, flags InputFlags)

@[c: 'igSetItemKeyOwner_Nil']
pub fn set_item_key_owner_nil(key Key)

@[c: 'igIsMouseDown_Nil']
pub fn is_mouse_down_nil(button MouseButton) bool

@[c: 'igIsMouseClicked_Bool']
pub fn is_mouse_clicked_bool(button MouseButton, repeat bool) bool

@[c: 'igIsMouseReleased_Nil']
pub fn is_mouse_released_nil(button MouseButton) bool

@[c: 'igIsMouseDoubleClicked_Nil']
pub fn is_mouse_double_clicked_nil(button MouseButton) bool

@[c: 'igIsMouseReleasedWithDelay']
pub fn is_mouse_released_with_delay(button MouseButton, delay f32) bool

@[c: 'igGetMouseClickedCount']
pub fn get_mouse_clicked_count(button MouseButton) int

@[c: 'igIsMouseHoveringRect']
pub fn is_mouse_hovering_rect(r_min ImVec2, r_max ImVec2, clip bool) bool

@[c: 'igIsMousePosValid']
pub fn is_mouse_pos_valid(mouse_pos &ImVec2) bool

@[c: 'igIsAnyMouseDown']
pub fn is_any_mouse_down() bool

@[c: 'igGetMousePos']
pub fn get_mouse_pos(p_out &ImVec2)

@[c: 'igGetMousePosOnOpeningCurrentPopup']
pub fn get_mouse_pos_on_opening_current_popup(p_out &ImVec2)

@[c: 'igIsMouseDragging']
pub fn is_mouse_dragging(button MouseButton, lock_threshold f32) bool

@[c: 'igGetMouseDragDelta']
pub fn get_mouse_drag_delta(p_out &ImVec2, button MouseButton, lock_threshold f32)

@[c: 'igResetMouseDragDelta']
pub fn reset_mouse_drag_delta(button MouseButton)

@[c: 'igGetMouseCursor']
pub fn get_mouse_cursor() MouseCursor

@[c: 'igSetMouseCursor']
pub fn set_mouse_cursor(cursor_type MouseCursor)

@[c: 'igSetNextFrameWantCaptureMouse']
pub fn set_next_frame_want_capture_mouse(want_capture_mouse bool)

@[c: 'igGetClipboardText']
pub fn get_clipboard_text() &i8

@[c: 'igSetClipboardText']
pub fn set_clipboard_text(text &i8)

@[c: 'igLoadIniSettingsFromDisk']
pub fn load_ini_settings_from_disk(ini_filename &i8)

@[c: 'igLoadIniSettingsFromMemory']
pub fn load_ini_settings_from_memory(ini_data &i8, ini_size usize)

@[c: 'igSaveIniSettingsToDisk']
pub fn save_ini_settings_to_disk(ini_filename &i8)

@[c: 'igSaveIniSettingsToMemory']
pub fn save_ini_settings_to_memory(out_ini_size &usize) &i8

@[c: 'igDebugTextEncoding']
pub fn debug_text_encoding(text &i8)

@[c: 'igDebugFlashStyleColor']
pub fn debug_flash_style_color(idx Col)

@[c: 'igDebugStartItemPicker']
pub fn debug_start_item_picker()

@[c: 'igDebugCheckVersionAndDataLayout']
pub fn debug_check_version_and_data_layout(version_str &i8, sz_io usize, sz_style usize, sz_vec2 usize, sz_vec4 usize, sz_drawvert usize, sz_drawidx usize) bool

@[c: 'igDebugLog']
@[c2v_variadic]
pub fn debug_log(fmt ...&i8)

@[c: 'igDebugLogV']
pub fn debug_log_v(fmt &i8, args Va_list)

@[c: 'igSetAllocatorFunctions']
pub fn set_allocator_functions(alloc_func MemAllocFunc, free_func MemFreeFunc, user_data voidptr)

@[c: 'igGetAllocatorFunctions']
pub fn get_allocator_functions(p_alloc_func &MemAllocFunc, p_free_func &MemFreeFunc, p_user_data &voidptr)

@[c: 'igMemAlloc']
pub fn mem_alloc(size usize) voidptr

@[c: 'igMemFree']
pub fn mem_free(ptr voidptr)

@[c: 'igUpdatePlatformWindows']
pub fn update_platform_windows()

@[c: 'igRenderPlatformWindowsDefault']
pub fn render_platform_windows_default(platform_render_arg voidptr, renderer_render_arg voidptr)

@[c: 'igDestroyPlatformWindows']
pub fn destroy_platform_windows()

@[c: 'igFindViewportByID']
pub fn find_viewport_by_id(id ID) &Viewport

@[c: 'igFindViewportByPlatformHandle']
pub fn find_viewport_by_platform_handle(platform_handle voidptr) &Viewport

@[c: 'TableSortSpecs_TableSortSpecs']
pub fn table_sort_specs_im_gui_table_sort_specs() &TableSortSpecs

@[c: 'TableSortSpecs_destroy']
pub fn table_sort_specs_destroy(self &TableSortSpecs)

@[c: 'TableColumnSortSpecs_TableColumnSortSpecs']
pub fn table_column_sort_specs_im_gui_table_column_sort_specs() &TableColumnSortSpecs

@[c: 'TableColumnSortSpecs_destroy']
pub fn table_column_sort_specs_destroy(self &TableColumnSortSpecs)

@[c: 'Style_Style']
pub fn style_im_gui_style() &Style

@[c: 'Style_destroy']
pub fn style_destroy(self &Style)

@[c: 'Style_ScaleAllSizes']
pub fn style_scale_all_sizes(self &Style, scale_factor f32)

@[c: 'IO_AddKeyEvent']
pub fn io_add_key_event(self &IO, key Key, down bool)

@[c: 'IO_AddKeyAnalogEvent']
pub fn io_add_key_analog_event(self &IO, key Key, down bool, v f32)

@[c: 'IO_AddMousePosEvent']
pub fn io_add_mouse_pos_event(self &IO, x f32, y f32)

@[c: 'IO_AddMouseButtonEvent']
pub fn io_add_mouse_button_event(self &IO, button int, down bool)

@[c: 'IO_AddMouseWheelEvent']
pub fn io_add_mouse_wheel_event(self &IO, wheel_x f32, wheel_y f32)

@[c: 'IO_AddMouseSourceEvent']
pub fn io_add_mouse_source_event(self &IO, source MouseSource)

@[c: 'IO_AddMouseViewportEvent']
pub fn io_add_mouse_viewport_event(self &IO, id ID)

@[c: 'IO_AddFocusEvent']
pub fn io_add_focus_event(self &IO, focused bool)

@[c: 'IO_AddInputCharacter']
pub fn io_add_input_character(self &IO, c u32)

@[c: 'IO_AddInputCharacterUTF16']
pub fn io_add_input_character_utf_16(self &IO, c ImWchar16)

@[c: 'IO_AddInputCharactersUTF8']
pub fn io_add_input_characters_utf_8(self &IO, str &i8)

@[c: 'IO_SetKeyEventNativeData']
pub fn io_set_key_event_native_data(self &IO, key Key, native_keycode int, native_scancode int, native_legacy_index int)

@[c: 'IO_SetAppAcceptingEvents']
pub fn io_set_app_accepting_events(self &IO, accepting_events bool)

@[c: 'IO_ClearEventsQueue']
pub fn io_clear_events_queue(self &IO)

@[c: 'IO_ClearInputKeys']
pub fn io_clear_input_keys(self &IO)

@[c: 'IO_ClearInputMouse']
pub fn io_clear_input_mouse(self &IO)

@[c: 'IO_IO']
pub fn io_im_gui_io() &IO

@[c: 'IO_destroy']
pub fn io_destroy(self &IO)

@[c: 'InputTextCallbackData_InputTextCallbackData']
pub fn input_text_callback_data_im_gui_input_text_callback_data() &InputTextCallbackData

@[c: 'InputTextCallbackData_destroy']
pub fn input_text_callback_data_destroy(self &InputTextCallbackData)

@[c: 'InputTextCallbackData_DeleteChars']
pub fn input_text_callback_data_delete_chars(self &InputTextCallbackData, pos int, bytes_count int)

@[c: 'InputTextCallbackData_InsertChars']
pub fn input_text_callback_data_insert_chars(self &InputTextCallbackData, pos int, text &i8, text_end &i8)

@[c: 'InputTextCallbackData_SelectAll']
pub fn input_text_callback_data_select_all(self &InputTextCallbackData)

@[c: 'InputTextCallbackData_ClearSelection']
pub fn input_text_callback_data_clear_selection(self &InputTextCallbackData)

@[c: 'InputTextCallbackData_HasSelection']
pub fn input_text_callback_data_has_selection(self &InputTextCallbackData) bool

@[c: 'WindowClass_WindowClass']
pub fn window_class_im_gui_window_class() &WindowClass

@[c: 'WindowClass_destroy']
pub fn window_class_destroy(self &WindowClass)

@[c: 'Payload_Payload']
pub fn payload_im_gui_payload() &Payload

@[c: 'Payload_destroy']
pub fn payload_destroy(self &Payload)

@[c: 'Payload_Clear']
pub fn payload_clear(self &Payload)

@[c: 'Payload_IsDataType']
pub fn payload_is_data_type(self &Payload, type_ &i8) bool

@[c: 'Payload_IsPreview']
pub fn payload_is_preview(self &Payload) bool

@[c: 'Payload_IsDelivery']
pub fn payload_is_delivery(self &Payload) bool

@[c: 'OnceUponAFrame_OnceUponAFrame']
pub fn once_upon_af_rame_im_gui_once_upon_af_rame() &OnceUponAFrame

@[c: 'OnceUponAFrame_destroy']
pub fn once_upon_af_rame_destroy(self &OnceUponAFrame)

@[c: 'TextFilter_TextFilter']
pub fn text_filter_im_gui_text_filter(default_filter &i8) &TextFilter

@[c: 'TextFilter_destroy']
pub fn text_filter_destroy(self &TextFilter)

@[c: 'TextFilter_Draw']
pub fn text_filter_draw(self &TextFilter, label &i8, width f32) bool

@[c: 'TextFilter_PassFilter']
pub fn text_filter_pass_filter(self &TextFilter, text &i8, text_end &i8) bool

@[c: 'TextFilter_Build']
pub fn text_filter_build(self &TextFilter)

@[c: 'TextFilter_Clear']
pub fn text_filter_clear(self &TextFilter)

@[c: 'TextFilter_IsActive']
pub fn text_filter_is_active(self &TextFilter) bool

@[c: 'TextRange_TextRange_Nil']
pub fn text_range_im_gui_text_range_nil() &TextRange

@[c: 'TextRange_destroy']
pub fn text_range_destroy(self &TextRange)

@[c: 'TextRange_TextRange_Str']
pub fn text_range_im_gui_text_range_str(_b &i8, _e &i8) &TextRange

@[c: 'TextRange_empty']
pub fn text_range_empty(self &TextRange) bool

@[c: 'TextRange_split']
pub fn text_range_split(self &TextRange, separator i8, out &ImVector_TextRange)

@[c: 'TextBuffer_TextBuffer']
pub fn text_buffer_im_gui_text_buffer() &TextBuffer

@[c: 'TextBuffer_destroy']
pub fn text_buffer_destroy(self &TextBuffer)

@[c: 'TextBuffer_begin']
pub fn text_buffer_begin(self &TextBuffer) &i8

@[c: 'TextBuffer_end']
pub fn text_buffer_end(self &TextBuffer) &i8

@[c: 'TextBuffer_size']
pub fn text_buffer_size(self &TextBuffer) int

@[c: 'TextBuffer_empty']
pub fn text_buffer_empty(self &TextBuffer) bool

@[c: 'TextBuffer_clear']
pub fn text_buffer_clear(self &TextBuffer)

@[c: 'TextBuffer_resize']
pub fn text_buffer_resize(self &TextBuffer, size int)

@[c: 'TextBuffer_reserve']
pub fn text_buffer_reserve(self &TextBuffer, capacity int)

@[c: 'TextBuffer_c_str']
pub fn text_buffer_c_str(self &TextBuffer) &i8

@[c: 'TextBuffer_append']
pub fn text_buffer_append(self &TextBuffer, str &i8, str_end &i8)

@[c: 'TextBuffer_appendfv']
pub fn text_buffer_appendfv(self &TextBuffer, fmt &i8, args Va_list)

@[c: 'StoragePair_StoragePair_Int']
pub fn storage_pair_im_gui_storage_pair_int(_key ID, _val int) &StoragePair

@[c: 'StoragePair_destroy']
pub fn storage_pair_destroy(self &StoragePair)

@[c: 'StoragePair_StoragePair_Float']
pub fn storage_pair_im_gui_storage_pair_float(_key ID, _val f32) &StoragePair

@[c: 'StoragePair_StoragePair_Ptr']
pub fn storage_pair_im_gui_storage_pair_ptr(_key ID, _val voidptr) &StoragePair

@[c: 'Storage_Clear']
pub fn storage_clear(self &Storage)

@[c: 'Storage_GetInt']
pub fn storage_get_int(self &Storage, key ID, default_val int) int

@[c: 'Storage_SetInt']
pub fn storage_set_int(self &Storage, key ID, val int)

@[c: 'Storage_GetBool']
pub fn storage_get_bool(self &Storage, key ID, default_val bool) bool

@[c: 'Storage_SetBool']
pub fn storage_set_bool(self &Storage, key ID, val bool)

@[c: 'Storage_GetFloat']
pub fn storage_get_float(self &Storage, key ID, default_val f32) f32

@[c: 'Storage_SetFloat']
pub fn storage_set_float(self &Storage, key ID, val f32)

@[c: 'Storage_GetVoidPtr']
pub fn storage_get_void_ptr(self &Storage, key ID) voidptr

@[c: 'Storage_SetVoidPtr']
pub fn storage_set_void_ptr(self &Storage, key ID, val voidptr)

@[c: 'Storage_GetIntRef']
pub fn storage_get_int_ref(self &Storage, key ID, default_val int) &int

@[c: 'Storage_GetBoolRef']
pub fn storage_get_bool_ref(self &Storage, key ID, default_val bool) &bool

@[c: 'Storage_GetFloatRef']
pub fn storage_get_float_ref(self &Storage, key ID, default_val f32) &f32

@[c: 'Storage_GetVoidPtrRef']
pub fn storage_get_void_ptr_ref(self &Storage, key ID, default_val voidptr) &voidptr

@[c: 'Storage_BuildSortByKey']
pub fn storage_build_sort_by_key(self &Storage)

@[c: 'Storage_SetAllInt']
pub fn storage_set_all_int(self &Storage, val int)

@[c: 'ListClipper_ListClipper']
pub fn list_clipper_im_gui_list_clipper() &ListClipper

@[c: 'ListClipper_destroy']
pub fn list_clipper_destroy(self &ListClipper)

@[c: 'ListClipper_Begin']
pub fn list_clipper_begin(self &ListClipper, items_count int, items_height f32)

@[c: 'ListClipper_End']
pub fn list_clipper_end(self &ListClipper)

@[c: 'ListClipper_Step']
pub fn list_clipper_step(self &ListClipper) bool

@[c: 'ListClipper_IncludeItemByIndex']
pub fn list_clipper_include_item_by_index(self &ListClipper, item_index int)

@[c: 'ListClipper_IncludeItemsByIndex']
pub fn list_clipper_include_items_by_index(self &ListClipper, item_begin int, item_end int)

@[c: 'ListClipper_SeekCursorForItem']
pub fn list_clipper_seek_cursor_for_item(self &ListClipper, item_index int)

@[c: 'ImColor_ImColor_Nil']
pub fn im_color_im_color_nil() &ImColor

@[c: 'ImColor_destroy']
pub fn im_color_destroy(self &ImColor)

@[c: 'ImColor_ImColor_Float']
pub fn im_color_im_color_float(r f32, g f32, b f32, a f32) &ImColor

@[c: 'ImColor_ImColor_Vec4']
pub fn im_color_im_color_vec4(col ImVec4) &ImColor

@[c: 'ImColor_ImColor_Int']
pub fn im_color_im_color_int(r int, g int, b int, a int) &ImColor

@[c: 'ImColor_ImColor_U32']
pub fn im_color_im_color_u32(rgba ImU32) &ImColor

@[c: 'ImColor_SetHSV']
pub fn im_color_set_hsv(self &ImColor, h f32, s f32, v f32, a f32)

@[c: 'ImColor_HSV']
pub fn im_color_hsv(p_out &ImColor, h f32, s f32, v f32, a f32)

@[c: 'SelectionBasicStorage_SelectionBasicStorage']
pub fn selection_basic_storage_im_gui_selection_basic_storage() &SelectionBasicStorage

@[c: 'SelectionBasicStorage_destroy']
pub fn selection_basic_storage_destroy(self &SelectionBasicStorage)

@[c: 'SelectionBasicStorage_ApplyRequests']
pub fn selection_basic_storage_apply_requests(self &SelectionBasicStorage, ms_io &MultiSelectIO)

@[c: 'SelectionBasicStorage_Contains']
pub fn selection_basic_storage_contains(self &SelectionBasicStorage, id ID) bool

@[c: 'SelectionBasicStorage_Clear']
pub fn selection_basic_storage_clear(self &SelectionBasicStorage)

@[c: 'SelectionBasicStorage_Swap']
pub fn selection_basic_storage_swap(self &SelectionBasicStorage, r &SelectionBasicStorage)

@[c: 'SelectionBasicStorage_SetItemSelected']
pub fn selection_basic_storage_set_item_selected(self &SelectionBasicStorage, id ID, selected bool)

@[c: 'SelectionBasicStorage_GetNextSelectedItem']
pub fn selection_basic_storage_get_next_selected_item(self &SelectionBasicStorage, opaque_it &voidptr, out_id &ID) bool

@[c: 'SelectionBasicStorage_GetStorageIdFromIndex']
pub fn selection_basic_storage_get_storage_id_from_index(self &SelectionBasicStorage, idx int) ID

@[c: 'SelectionExternalStorage_SelectionExternalStorage']
pub fn selection_external_storage_im_gui_selection_external_storage() &SelectionExternalStorage

@[c: 'SelectionExternalStorage_destroy']
pub fn selection_external_storage_destroy(self &SelectionExternalStorage)

@[c: 'SelectionExternalStorage_ApplyRequests']
pub fn selection_external_storage_apply_requests(self &SelectionExternalStorage, ms_io &MultiSelectIO)

@[c: 'ImDrawCmd_ImDrawCmd']
pub fn im_draw_cmd_im_draw_cmd() &ImDrawCmd

@[c: 'ImDrawCmd_destroy']
pub fn im_draw_cmd_destroy(self &ImDrawCmd)

@[c: 'ImDrawCmd_GetTexID']
pub fn im_draw_cmd_get_tex_id(self &ImDrawCmd) ImTextureID

@[c: 'ImDrawListSplitter_ImDrawListSplitter']
pub fn im_draw_list_splitter_im_draw_list_splitter() &ImDrawListSplitter

@[c: 'ImDrawListSplitter_destroy']
pub fn im_draw_list_splitter_destroy(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_Clear']
pub fn im_draw_list_splitter_clear(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_ClearFreeMemory']
pub fn im_draw_list_splitter_clear_free_memory(self &ImDrawListSplitter)

@[c: 'ImDrawListSplitter_Split']
pub fn im_draw_list_splitter_split(self &ImDrawListSplitter, draw_list &ImDrawList, count int)

@[c: 'ImDrawListSplitter_Merge']
pub fn im_draw_list_splitter_merge(self &ImDrawListSplitter, draw_list &ImDrawList)

@[c: 'ImDrawListSplitter_SetCurrentChannel']
pub fn im_draw_list_splitter_set_current_channel(self &ImDrawListSplitter, draw_list &ImDrawList, channel_idx int)

@[c: 'ImDrawList_ImDrawList']
pub fn im_draw_list_im_draw_list(shared_data &ImDrawListSharedData) &ImDrawList

@[c: 'ImDrawList_destroy']
pub fn im_draw_list_destroy(self &ImDrawList)

@[c: 'ImDrawList_PushClipRect']
pub fn im_draw_list_push_clip_rect(self &ImDrawList, clip_rect_min ImVec2, clip_rect_max ImVec2, intersect_with_current_clip_rect bool)

@[c: 'ImDrawList_PushClipRectFullScreen']
pub fn im_draw_list_push_clip_rect_full_screen(self &ImDrawList)

@[c: 'ImDrawList_PopClipRect']
pub fn im_draw_list_pop_clip_rect(self &ImDrawList)

@[c: 'ImDrawList_PushTextureID']
pub fn im_draw_list_push_texture_id(self &ImDrawList, texture_id ImTextureID)

@[c: 'ImDrawList_PopTextureID']
pub fn im_draw_list_pop_texture_id(self &ImDrawList)

@[c: 'ImDrawList_GetClipRectMin']
pub fn im_draw_list_get_clip_rect_min(p_out &ImVec2, self &ImDrawList)

@[c: 'ImDrawList_GetClipRectMax']
pub fn im_draw_list_get_clip_rect_max(p_out &ImVec2, self &ImDrawList)

@[c: 'ImDrawList_AddLine']
pub fn im_draw_list_add_line(self &ImDrawList, p1 ImVec2, p2 ImVec2, col ImU32, thickness f32)

@[c: 'ImDrawList_AddRect']
pub fn im_draw_list_add_rect(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags, thickness f32)

@[c: 'ImDrawList_AddRectFilled']
pub fn im_draw_list_add_rect_filled(self &ImDrawList, p_min ImVec2, p_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags)

@[c: 'ImDrawList_AddRectFilledMultiColor']
pub fn im_draw_list_add_rect_filled_multi_color(self &ImDrawList, p_min ImVec2, p_max ImVec2, col_upr_left ImU32, col_upr_right ImU32, col_bot_right ImU32, col_bot_left ImU32)

@[c: 'ImDrawList_AddQuad']
pub fn im_draw_list_add_quad(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32, thickness f32)

@[c: 'ImDrawList_AddQuadFilled']
pub fn im_draw_list_add_quad_filled(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32)

@[c: 'ImDrawList_AddTriangle']
pub fn im_draw_list_add_triangle(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32, thickness f32)

@[c: 'ImDrawList_AddTriangleFilled']
pub fn im_draw_list_add_triangle_filled(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32)

@[c: 'ImDrawList_AddCircle']
pub fn im_draw_list_add_circle(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int, thickness f32)

@[c: 'ImDrawList_AddCircleFilled']
pub fn im_draw_list_add_circle_filled(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

@[c: 'ImDrawList_AddNgon']
pub fn im_draw_list_add_ngon(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int, thickness f32)

@[c: 'ImDrawList_AddNgonFilled']
pub fn im_draw_list_add_ngon_filled(self &ImDrawList, center ImVec2, radius f32, col ImU32, num_segments int)

@[c: 'ImDrawList_AddEllipse']
pub fn im_draw_list_add_ellipse(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32, rot f32, num_segments int, thickness f32)

@[c: 'ImDrawList_AddEllipseFilled']
pub fn im_draw_list_add_ellipse_filled(self &ImDrawList, center ImVec2, radius ImVec2, col ImU32, rot f32, num_segments int)

@[c: 'ImDrawList_AddText_Vec2']
pub fn im_draw_list_add_text_vec2(self &ImDrawList, pos ImVec2, col ImU32, text_begin &i8, text_end &i8)

@[c: 'ImDrawList_AddText_FontPtr']
pub fn im_draw_list_add_text_font_ptr(self &ImDrawList, font &ImFont, font_size f32, pos ImVec2, col ImU32, text_begin &i8, text_end &i8, wrap_width f32, cpu_fine_clip_rect &ImVec4)

@[c: 'ImDrawList_AddBezierCubic']
pub fn im_draw_list_add_bezier_cubic(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, col ImU32, thickness f32, num_segments int)

@[c: 'ImDrawList_AddBezierQuadratic']
pub fn im_draw_list_add_bezier_quadratic(self &ImDrawList, p1 ImVec2, p2 ImVec2, p3 ImVec2, col ImU32, thickness f32, num_segments int)

@[c: 'ImDrawList_AddPolyline']
pub fn im_draw_list_add_polyline(self &ImDrawList, points &ImVec2, num_points int, col ImU32, flags ImDrawFlags, thickness f32)

@[c: 'ImDrawList_AddConvexPolyFilled']
pub fn im_draw_list_add_convex_poly_filled(self &ImDrawList, points &ImVec2, num_points int, col ImU32)

@[c: 'ImDrawList_AddConcavePolyFilled']
pub fn im_draw_list_add_concave_poly_filled(self &ImDrawList, points &ImVec2, num_points int, col ImU32)

@[c: 'ImDrawList_AddImage']
pub fn im_draw_list_add_image(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2, uv_min ImVec2, uv_max ImVec2, col ImU32)

@[c: 'ImDrawList_AddImageQuad']
pub fn im_draw_list_add_image_quad(self &ImDrawList, user_texture_id ImTextureID, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, uv1 ImVec2, uv2 ImVec2, uv3 ImVec2, uv4 ImVec2, col ImU32)

@[c: 'ImDrawList_AddImageRounded']
pub fn im_draw_list_add_image_rounded(self &ImDrawList, user_texture_id ImTextureID, p_min ImVec2, p_max ImVec2, uv_min ImVec2, uv_max ImVec2, col ImU32, rounding f32, flags ImDrawFlags)

@[c: 'ImDrawList_PathClear']
pub fn im_draw_list_path_clear(self &ImDrawList)

@[c: 'ImDrawList_PathLineTo']
pub fn im_draw_list_path_line_to(self &ImDrawList, pos ImVec2)

@[c: 'ImDrawList_PathLineToMergeDuplicate']
pub fn im_draw_list_path_line_to_merge_duplicate(self &ImDrawList, pos ImVec2)

@[c: 'ImDrawList_PathFillConvex']
pub fn im_draw_list_path_fill_convex(self &ImDrawList, col ImU32)

@[c: 'ImDrawList_PathFillConcave']
pub fn im_draw_list_path_fill_concave(self &ImDrawList, col ImU32)

@[c: 'ImDrawList_PathStroke']
pub fn im_draw_list_path_stroke(self &ImDrawList, col ImU32, flags ImDrawFlags, thickness f32)

@[c: 'ImDrawList_PathArcTo']
pub fn im_draw_list_path_arc_to(self &ImDrawList, center ImVec2, radius f32, a_min f32, a_max f32, num_segments int)

@[c: 'ImDrawList_PathArcToFast']
pub fn im_draw_list_path_arc_to_fast(self &ImDrawList, center ImVec2, radius f32, a_min_of_12 int, a_max_of_12 int)

@[c: 'ImDrawList_PathEllipticalArcTo']
pub fn im_draw_list_path_elliptical_arc_to(self &ImDrawList, center ImVec2, radius ImVec2, rot f32, a_min f32, a_max f32, num_segments int)

@[c: 'ImDrawList_PathBezierCubicCurveTo']
pub fn im_draw_list_path_bezier_cubic_curve_to(self &ImDrawList, p2 ImVec2, p3 ImVec2, p4 ImVec2, num_segments int)

@[c: 'ImDrawList_PathBezierQuadraticCurveTo']
pub fn im_draw_list_path_bezier_quadratic_curve_to(self &ImDrawList, p2 ImVec2, p3 ImVec2, num_segments int)

@[c: 'ImDrawList_PathRect']
pub fn im_draw_list_path_rect(self &ImDrawList, rect_min ImVec2, rect_max ImVec2, rounding f32, flags ImDrawFlags)

@[c: 'ImDrawList_AddCallback']
pub fn im_draw_list_add_callback(self &ImDrawList, callback ImDrawCallback, userdata voidptr, userdata_size usize)

@[c: 'ImDrawList_AddDrawCmd']
pub fn im_draw_list_add_draw_cmd(self &ImDrawList)

@[c: 'ImDrawList_CloneOutput']
pub fn im_draw_list_clone_output(self &ImDrawList) &ImDrawList

@[c: 'ImDrawList_ChannelsSplit']
pub fn im_draw_list_channels_split(self &ImDrawList, count int)

@[c: 'ImDrawList_ChannelsMerge']
pub fn im_draw_list_channels_merge(self &ImDrawList)

@[c: 'ImDrawList_ChannelsSetCurrent']
pub fn im_draw_list_channels_set_current(self &ImDrawList, n int)

@[c: 'ImDrawList_PrimReserve']
pub fn im_draw_list_prim_reserve(self &ImDrawList, idx_count int, vtx_count int)

@[c: 'ImDrawList_PrimUnreserve']
pub fn im_draw_list_prim_unreserve(self &ImDrawList, idx_count int, vtx_count int)

@[c: 'ImDrawList_PrimRect']
pub fn im_draw_list_prim_rect(self &ImDrawList, a ImVec2, b ImVec2, col ImU32)

@[c: 'ImDrawList_PrimRectUV']
pub fn im_draw_list_prim_rect_uv(self &ImDrawList, a ImVec2, b ImVec2, uv_a ImVec2, uv_b ImVec2, col ImU32)

@[c: 'ImDrawList_PrimQuadUV']
pub fn im_draw_list_prim_quad_uv(self &ImDrawList, a ImVec2, b ImVec2, c ImVec2, d ImVec2, uv_a ImVec2, uv_b ImVec2, uv_c ImVec2, uv_d ImVec2, col ImU32)

@[c: 'ImDrawList_PrimWriteVtx']
pub fn im_draw_list_prim_write_vtx(self &ImDrawList, pos ImVec2, uv ImVec2, col ImU32)

@[c: 'ImDrawList_PrimWriteIdx']
pub fn im_draw_list_prim_write_idx(self &ImDrawList, idx ImDrawIdx)

@[c: 'ImDrawList_PrimVtx']
pub fn im_draw_list_prim_vtx(self &ImDrawList, pos ImVec2, uv ImVec2, col ImU32)

@[c: 'ImDrawList__ResetForNewFrame']
pub fn im_draw_list__reset_for_new_frame(self &ImDrawList)

@[c: 'ImDrawList__ClearFreeMemory']
pub fn im_draw_list__clear_free_memory(self &ImDrawList)

@[c: 'ImDrawList__PopUnusedDrawCmd']
pub fn im_draw_list__pop_unused_draw_cmd(self &ImDrawList)

@[c: 'ImDrawList__TryMergeDrawCmds']
pub fn im_draw_list__try_merge_draw_cmds(self &ImDrawList)

@[c: 'ImDrawList__OnChangedClipRect']
pub fn im_draw_list__on_changed_clip_rect(self &ImDrawList)

@[c: 'ImDrawList__OnChangedTextureID']
pub fn im_draw_list__on_changed_texture_id(self &ImDrawList)

@[c: 'ImDrawList__OnChangedVtxOffset']
pub fn im_draw_list__on_changed_vtx_offset(self &ImDrawList)

@[c: 'ImDrawList__SetTextureID']
pub fn im_draw_list__set_texture_id(self &ImDrawList, texture_id ImTextureID)

@[c: 'ImDrawList__CalcCircleAutoSegmentCount']
pub fn im_draw_list__calc_circle_auto_segment_count(self &ImDrawList, radius f32) int

@[c: 'ImDrawList__PathArcToFastEx']
pub fn im_draw_list__path_arc_to_fast_ex(self &ImDrawList, center ImVec2, radius f32, a_min_sample int, a_max_sample int, a_step int)

@[c: 'ImDrawList__PathArcToN']
pub fn im_draw_list__path_arc_to_n(self &ImDrawList, center ImVec2, radius f32, a_min f32, a_max f32, num_segments int)

@[c: 'ImDrawData_ImDrawData']
pub fn im_draw_data_im_draw_data() &ImDrawData

@[c: 'ImDrawData_destroy']
pub fn im_draw_data_destroy(self &ImDrawData)

@[c: 'ImDrawData_Clear']
pub fn im_draw_data_clear(self &ImDrawData)

@[c: 'ImDrawData_AddDrawList']
pub fn im_draw_data_add_draw_list(self &ImDrawData, draw_list &ImDrawList)

@[c: 'ImDrawData_DeIndexAllBuffers']
pub fn im_draw_data_de_index_all_buffers(self &ImDrawData)

@[c: 'ImDrawData_ScaleClipRects']
pub fn im_draw_data_scale_clip_rects(self &ImDrawData, fb_scale ImVec2)

@[c: 'ImFontConfig_ImFontConfig']
pub fn im_font_config_im_font_config() &ImFontConfig

@[c: 'ImFontConfig_destroy']
pub fn im_font_config_destroy(self &ImFontConfig)

@[c: 'ImFontGlyphRangesBuilder_ImFontGlyphRangesBuilder']
pub fn im_font_glyph_ranges_builder_im_font_glyph_ranges_builder() &ImFontGlyphRangesBuilder

@[c: 'ImFontGlyphRangesBuilder_destroy']
pub fn im_font_glyph_ranges_builder_destroy(self &ImFontGlyphRangesBuilder)

@[c: 'ImFontGlyphRangesBuilder_Clear']
pub fn im_font_glyph_ranges_builder_clear(self &ImFontGlyphRangesBuilder)

@[c: 'ImFontGlyphRangesBuilder_GetBit']
pub fn im_font_glyph_ranges_builder_get_bit(self &ImFontGlyphRangesBuilder, n usize) bool

@[c: 'ImFontGlyphRangesBuilder_SetBit']
pub fn im_font_glyph_ranges_builder_set_bit(self &ImFontGlyphRangesBuilder, n usize)

@[c: 'ImFontGlyphRangesBuilder_AddChar']
pub fn im_font_glyph_ranges_builder_add_char(self &ImFontGlyphRangesBuilder, c ImWchar)

@[c: 'ImFontGlyphRangesBuilder_AddText']
pub fn im_font_glyph_ranges_builder_add_text(self &ImFontGlyphRangesBuilder, text &i8, text_end &i8)

@[c: 'ImFontGlyphRangesBuilder_AddRanges']
pub fn im_font_glyph_ranges_builder_add_ranges(self &ImFontGlyphRangesBuilder, ranges &ImWchar)

@[c: 'ImFontGlyphRangesBuilder_BuildRanges']
pub fn im_font_glyph_ranges_builder_build_ranges(self &ImFontGlyphRangesBuilder, out_ranges &ImVector_ImWchar)

@[c: 'ImFontAtlasCustomRect_ImFontAtlasCustomRect']
pub fn im_font_atlas_custom_rect_im_font_atlas_custom_rect() &ImFontAtlasCustomRect

@[c: 'ImFontAtlasCustomRect_destroy']
pub fn im_font_atlas_custom_rect_destroy(self &ImFontAtlasCustomRect)

@[c: 'ImFontAtlasCustomRect_IsPacked']
pub fn im_font_atlas_custom_rect_is_packed(self &ImFontAtlasCustomRect) bool

@[c: 'ImFontAtlas_ImFontAtlas']
pub fn im_font_atlas_im_font_atlas() &ImFontAtlas

@[c: 'ImFontAtlas_destroy']
pub fn im_font_atlas_destroy(self &ImFontAtlas)

@[c: 'ImFontAtlas_AddFont']
pub fn im_font_atlas_add_font(self &ImFontAtlas, font_cfg &ImFontConfig) &ImFont

@[c: 'ImFontAtlas_AddFontDefault']
pub fn im_font_atlas_add_font_default(self &ImFontAtlas, font_cfg &ImFontConfig) &ImFont

@[c: 'ImFontAtlas_AddFontFromFileTTF']
pub fn im_font_atlas_add_font_from_file_ttf(self &ImFontAtlas, filename &i8, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &ImWchar) &ImFont

@[c: 'ImFontAtlas_AddFontFromMemoryTTF']
pub fn im_font_atlas_add_font_from_memory_ttf(self &ImFontAtlas, font_data voidptr, font_data_size int, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &ImWchar) &ImFont

@[c: 'ImFontAtlas_AddFontFromMemoryCompressedTTF']
pub fn im_font_atlas_add_font_from_memory_compressed_ttf(self &ImFontAtlas, compressed_font_data voidptr, compressed_font_data_size int, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &ImWchar) &ImFont

@[c: 'ImFontAtlas_AddFontFromMemoryCompressedBase85TTF']
pub fn im_font_atlas_add_font_from_memory_compressed_base85_ttf(self &ImFontAtlas, compressed_font_data_base85 &i8, size_pixels f32, font_cfg &ImFontConfig, glyph_ranges &ImWchar) &ImFont

@[c: 'ImFontAtlas_ClearInputData']
pub fn im_font_atlas_clear_input_data(self &ImFontAtlas)

@[c: 'ImFontAtlas_ClearFonts']
pub fn im_font_atlas_clear_fonts(self &ImFontAtlas)

@[c: 'ImFontAtlas_ClearTexData']
pub fn im_font_atlas_clear_tex_data(self &ImFontAtlas)

@[c: 'ImFontAtlas_Clear']
pub fn im_font_atlas_clear(self &ImFontAtlas)

@[c: 'ImFontAtlas_Build']
pub fn im_font_atlas_build(self &ImFontAtlas) bool

@[c: 'ImFontAtlas_GetTexDataAsAlpha8']
pub fn im_font_atlas_get_tex_data_as_alpha8(self &ImFontAtlas, out_pixels &&u8, out_width &int, out_height &int, out_bytes_per_pixel &int)

@[c: 'ImFontAtlas_GetTexDataAsRGBA32']
pub fn im_font_atlas_get_tex_data_as_rgba_32(self &ImFontAtlas, out_pixels &&u8, out_width &int, out_height &int, out_bytes_per_pixel &int)

@[c: 'ImFontAtlas_IsBuilt']
pub fn im_font_atlas_is_built(self &ImFontAtlas) bool

@[c: 'ImFontAtlas_SetTexID']
pub fn im_font_atlas_set_tex_id(self &ImFontAtlas, id ImTextureID)

@[c: 'ImFontAtlas_GetGlyphRangesDefault']
pub fn im_font_atlas_get_glyph_ranges_default(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesGreek']
pub fn im_font_atlas_get_glyph_ranges_greek(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesKorean']
pub fn im_font_atlas_get_glyph_ranges_korean(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesJapanese']
pub fn im_font_atlas_get_glyph_ranges_japanese(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesChineseFull']
pub fn im_font_atlas_get_glyph_ranges_chinese_full(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesChineseSimplifiedCommon']
pub fn im_font_atlas_get_glyph_ranges_chinese_simplified_common(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesCyrillic']
pub fn im_font_atlas_get_glyph_ranges_cyrillic(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesThai']
pub fn im_font_atlas_get_glyph_ranges_thai(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_GetGlyphRangesVietnamese']
pub fn im_font_atlas_get_glyph_ranges_vietnamese(self &ImFontAtlas) &ImWchar

@[c: 'ImFontAtlas_AddCustomRectRegular']
pub fn im_font_atlas_add_custom_rect_regular(self &ImFontAtlas, width int, height int) int

@[c: 'ImFontAtlas_AddCustomRectFontGlyph']
pub fn im_font_atlas_add_custom_rect_font_glyph(self &ImFontAtlas, font &ImFont, id ImWchar, width int, height int, advance_x f32, offset ImVec2) int

@[c: 'ImFontAtlas_GetCustomRectByIndex']
pub fn im_font_atlas_get_custom_rect_by_index(self &ImFontAtlas, index int) &ImFontAtlasCustomRect

@[c: 'ImFontAtlas_CalcCustomRectUV']
pub fn im_font_atlas_calc_custom_rect_uv(self &ImFontAtlas, rect &ImFontAtlasCustomRect, out_uv_min &ImVec2, out_uv_max &ImVec2)

@[c: 'ImFont_ImFont']
pub fn im_font_im_font() &ImFont

@[c: 'ImFont_destroy']
pub fn im_font_destroy(self &ImFont)

@[c: 'ImFont_FindGlyph']
pub fn im_font_find_glyph(self &ImFont, c ImWchar) &ImFontGlyph

@[c: 'ImFont_FindGlyphNoFallback']
pub fn im_font_find_glyph_no_fallback(self &ImFont, c ImWchar) &ImFontGlyph

@[c: 'ImFont_GetCharAdvance']
pub fn im_font_get_char_advance(self &ImFont, c ImWchar) f32

@[c: 'ImFont_IsLoaded']
pub fn im_font_is_loaded(self &ImFont) bool

@[c: 'ImFont_GetDebugName']
pub fn im_font_get_debug_name(self &ImFont) &i8

@[c: 'ImFont_CalcTextSizeA']
pub fn im_font_calc_text_size_a(p_out &ImVec2, self &ImFont, size f32, max_width f32, wrap_width f32, text_begin &i8, text_end &i8, remaining &&u8)

@[c: 'ImFont_CalcWordWrapPositionA']
pub fn im_font_calc_word_wrap_position_a(self &ImFont, scale f32, text &i8, text_end &i8, wrap_width f32) &i8

@[c: 'ImFont_RenderChar']
pub fn im_font_render_char(self &ImFont, draw_list &ImDrawList, size f32, pos ImVec2, col ImU32, c ImWchar)

@[c: 'ImFont_RenderText']
pub fn im_font_render_text(self &ImFont, draw_list &ImDrawList, size f32, pos ImVec2, col ImU32, clip_rect ImVec4, text_begin &i8, text_end &i8, wrap_width f32, cpu_fine_clip bool)

@[c: 'ImFont_BuildLookupTable']
pub fn im_font_build_lookup_table(self &ImFont)

@[c: 'ImFont_ClearOutputData']
pub fn im_font_clear_output_data(self &ImFont)

@[c: 'ImFont_GrowIndex']
pub fn im_font_grow_index(self &ImFont, new_size int)

@[c: 'ImFont_AddGlyph']
pub fn im_font_add_glyph(self &ImFont, src_cfg &ImFontConfig, c ImWchar, x0 f32, y0 f32, x1 f32, y1 f32, u0 f32, v0 f32, u1 f32, v1 f32, advance_x f32)

@[c: 'ImFont_AddRemapChar']
pub fn im_font_add_remap_char(self &ImFont, dst ImWchar, src ImWchar, overwrite_dst bool)

@[c: 'ImFont_IsGlyphRangeUnused']
pub fn im_font_is_glyph_range_unused(self &ImFont, c_begin u32, c_last u32) bool

@[c: 'Viewport_Viewport']
pub fn viewport_im_gui_viewport() &Viewport

@[c: 'Viewport_destroy']
pub fn viewport_destroy(self &Viewport)

@[c: 'Viewport_GetCenter']
pub fn viewport_get_center(p_out &ImVec2, self &Viewport)

@[c: 'Viewport_GetWorkCenter']
pub fn viewport_get_work_center(p_out &ImVec2, self &Viewport)

@[c: 'PlatformIO_PlatformIO']
pub fn platform_io_im_gui_platform_io() &PlatformIO

@[c: 'PlatformIO_destroy']
pub fn platform_io_destroy(self &PlatformIO)

@[c: 'PlatformMonitor_PlatformMonitor']
pub fn platform_monitor_im_gui_platform_monitor() &PlatformMonitor

@[c: 'PlatformMonitor_destroy']
pub fn platform_monitor_destroy(self &PlatformMonitor)

@[c: 'PlatformImeData_PlatformImeData']
pub fn platform_ime_data_im_gui_platform_ime_data() &PlatformImeData

@[c: 'PlatformImeData_destroy']
pub fn platform_ime_data_destroy(self &PlatformImeData)

@[c: 'igImHashData']
pub fn im_hash_data(data voidptr, data_size usize, seed ID) ID

@[c: 'igImHashStr']
pub fn im_hash_str(data &i8, data_size usize, seed ID) ID

@[c: 'igImQsort']
pub fn im_qsort(base voidptr, count usize, size_of_element usize, compare_func fn (voidptr, voidptr) int)

@[c: 'igImAlphaBlendColors']
pub fn im_alpha_blend_colors(col_a ImU32, col_b ImU32) ImU32

@[c: 'igImIsPowerOfTwo_Int']
pub fn im_is_power_of_two_int(v int) bool

@[c: 'igImIsPowerOfTwo_U64']
pub fn im_is_power_of_two_u64(v ImU64) bool

@[c: 'igImUpperPowerOfTwo']
pub fn im_upper_power_of_two(v int) int

@[c: 'igImCountSetBits']
pub fn im_count_set_bits(v u32) u32

@[c: 'igImStricmp']
pub fn im_stricmp(str1 &i8, str2 &i8) int

@[c: 'igImStrnicmp']
pub fn im_strnicmp(str1 &i8, str2 &i8, count usize) int

@[c: 'igImStrncpy']
pub fn im_strncpy(dst &i8, src &i8, count usize)

@[c: 'igImStrdup']
pub fn im_strdup(str &i8) &i8

@[c: 'igImStrdupcpy']
pub fn im_strdupcpy(dst &i8, p_dst_size &usize, str &i8) &i8

@[c: 'igImStrchrRange']
pub fn im_strchr_range(str_begin &i8, str_end &i8, c i8) &i8

@[c: 'igImStreolRange']
pub fn im_streol_range(str &i8, str_end &i8) &i8

@[c: 'igImStristr']
pub fn im_stristr(haystack &i8, haystack_end &i8, needle &i8, needle_end &i8) &i8

@[c: 'igImStrTrimBlanks']
pub fn im_str_trim_blanks(str &i8)

@[c: 'igImStrSkipBlank']
pub fn im_str_skip_blank(str &i8) &i8

@[c: 'igImStrlenW']
pub fn im_strlen_w(str &ImWchar) int

@[c: 'igImStrbol']
pub fn im_strbol(buf_mid_line &i8, buf_begin &i8) &i8

@[c: 'igImToUpper']
pub fn im_to_upper(c i8) i8

@[c: 'igImCharIsBlankA']
pub fn im_char_is_blank_a(c i8) bool

@[c: 'igImCharIsBlankW']
pub fn im_char_is_blank_w(c u32) bool

@[c: 'igImCharIsXdigitA']
pub fn im_char_is_xdigit_a(c i8) bool

@[c: 'igImFormatString']
@[c2v_variadic]
pub fn im_format_string(buf &i8, buf_size usize, fmt ...&i8) int

@[c: 'igImFormatStringV']
pub fn im_format_string_v(buf &i8, buf_size usize, fmt &i8, args Va_list) int

@[c: 'igImFormatStringToTempBuffer']
@[c2v_variadic]
pub fn im_format_string_to_temp_buffer(out_buf &&u8, out_buf_end &&u8, fmt ...&i8)

@[c: 'igImFormatStringToTempBufferV']
pub fn im_format_string_to_temp_buffer_v(out_buf &&u8, out_buf_end &&u8, fmt &i8, args Va_list)

@[c: 'igImParseFormatFindStart']
pub fn im_parse_format_find_start(format &i8) &i8

@[c: 'igImParseFormatFindEnd']
pub fn im_parse_format_find_end(format &i8) &i8

@[c: 'igImParseFormatTrimDecorations']
pub fn im_parse_format_trim_decorations(format &i8, buf &i8, buf_size usize) &i8

@[c: 'igImParseFormatSanitizeForPrinting']
pub fn im_parse_format_sanitize_for_printing(fmt_in &i8, fmt_out &i8, fmt_out_size usize)

@[c: 'igImParseFormatSanitizeForScanning']
pub fn im_parse_format_sanitize_for_scanning(fmt_in &i8, fmt_out &i8, fmt_out_size usize) &i8

@[c: 'igImParseFormatPrecision']
pub fn im_parse_format_precision(format &i8, default_value int) int

@[c: 'igImTextCharToUtf8']
pub fn im_text_char_to_utf8(out_buf &i8, c u32) &i8

@[c: 'igImTextStrToUtf8']
pub fn im_text_str_to_utf8(out_buf &i8, out_buf_size int, in_text &ImWchar, in_text_end &ImWchar) int

@[c: 'igImTextCharFromUtf8']
pub fn im_text_char_from_utf8(out_char &u32, in_text &i8, in_text_end &i8) int

@[c: 'igImTextStrFromUtf8']
pub fn im_text_str_from_utf8(out_buf &ImWchar, out_buf_size int, in_text &i8, in_text_end &i8, in_remaining &&u8) int

@[c: 'igImTextCountCharsFromUtf8']
pub fn im_text_count_chars_from_utf8(in_text &i8, in_text_end &i8) int

@[c: 'igImTextCountUtf8BytesFromChar']
pub fn im_text_count_utf8_bytes_from_char(in_text &i8, in_text_end &i8) int

@[c: 'igImTextCountUtf8BytesFromStr']
pub fn im_text_count_utf8_bytes_from_str(in_text &ImWchar, in_text_end &ImWchar) int

@[c: 'igImTextFindPreviousUtf8Codepoint']
pub fn im_text_find_previous_utf8_codepoint(in_text_start &i8, in_text_curr &i8) &i8

@[c: 'igImTextCountLines']
pub fn im_text_count_lines(in_text &i8, in_text_end &i8) int

@[c: 'igImFileOpen']
pub fn im_file_open(filename &i8, mode &i8) ImFileHandle

@[c: 'igImFileClose']
pub fn im_file_close(file ImFileHandle) bool

@[c: 'igImFileGetSize']
pub fn im_file_get_size(file ImFileHandle) ImU64

@[c: 'igImFileRead']
pub fn im_file_read(data voidptr, size ImU64, count ImU64, file ImFileHandle) ImU64

@[c: 'igImFileWrite']
pub fn im_file_write(data voidptr, size ImU64, count ImU64, file ImFileHandle) ImU64

@[c: 'igImFileLoadToMemory']
pub fn im_file_load_to_memory(filename &i8, mode &i8, out_file_size &usize, padding_bytes int) voidptr

@[c: 'igImPow_Float']
pub fn im_pow_float(x f32, y f32) f32

@[c: 'igImPow_double']
pub fn im_pow_double(x f64, y f64) f64

@[c: 'igImLog_Float']
pub fn im_log_float(x f32) f32

@[c: 'igImLog_double']
pub fn im_log_double(x f64) f64

@[c: 'igImAbs_Int']
pub fn im_abs_int(x int) int

@[c: 'igImAbs_Float']
pub fn im_abs_float(x f32) f32

@[c: 'igImAbs_double']
pub fn im_abs_double(x f64) f64

@[c: 'igImSign_Float']
pub fn im_sign_float(x f32) f32

@[c: 'igImSign_double']
pub fn im_sign_double(x f64) f64

@[c: 'igImRsqrt_Float']
pub fn im_rsqrt_float(x f32) f32

@[c: 'igImRsqrt_double']
pub fn im_rsqrt_double(x f64) f64

@[c: 'igImMin']
pub fn im_min(p_out &ImVec2, lhs ImVec2, rhs ImVec2)

@[c: 'igImMax']
pub fn im_max(p_out &ImVec2, lhs ImVec2, rhs ImVec2)

@[c: 'igImClamp']
pub fn im_clamp(p_out &ImVec2, v ImVec2, mn ImVec2, mx ImVec2)

@[c: 'igImLerp_Vec2Float']
pub fn im_lerp_vec2_float(p_out &ImVec2, a ImVec2, b ImVec2, t f32)

@[c: 'igImLerp_Vec2Vec2']
pub fn im_lerp_vec2_vec2(p_out &ImVec2, a ImVec2, b ImVec2, t ImVec2)

@[c: 'igImLerp_Vec4']
pub fn im_lerp_vec4(p_out &ImVec4, a ImVec4, b ImVec4, t f32)

@[c: 'igImSaturate']
pub fn im_saturate(f f32) f32

@[c: 'igImLengthSqr_Vec2']
pub fn im_length_sqr_vec2(lhs ImVec2) f32

@[c: 'igImLengthSqr_Vec4']
pub fn im_length_sqr_vec4(lhs ImVec4) f32

@[c: 'igImInvLength']
pub fn im_inv_length(lhs ImVec2, fail_value f32) f32

@[c: 'igImTrunc_Float']
pub fn im_trunc_float(f f32) f32

@[c: 'igImTrunc_Vec2']
pub fn im_trunc_vec2(p_out &ImVec2, v ImVec2)

@[c: 'igImFloor_Float']
pub fn im_floor_float(f f32) f32

@[c: 'igImFloor_Vec2']
pub fn im_floor_vec2(p_out &ImVec2, v ImVec2)

@[c: 'igImModPositive']
pub fn im_mod_positive(a int, b int) int

@[c: 'igImDot']
pub fn im_dot(a ImVec2, b ImVec2) f32

@[c: 'igImRotate']
pub fn im_rotate(p_out &ImVec2, v ImVec2, cos_a f32, sin_a f32)

@[c: 'igImLinearSweep']
pub fn im_linear_sweep(current f32, target f32, speed f32) f32

@[c: 'igImLinearRemapClamp']
pub fn im_linear_remap_clamp(s0 f32, s1 f32, d0 f32, d1 f32, x f32) f32

@[c: 'igImMul']
pub fn im_mul(p_out &ImVec2, lhs ImVec2, rhs ImVec2)

@[c: 'igImIsFloatAboveGuaranteedIntegerPrecision']
pub fn im_is_float_above_guaranteed_integer_precision(f f32) bool

@[c: 'igImExponentialMovingAverage']
pub fn im_exponential_moving_average(avg f32, sample f32, n int) f32

@[c: 'igImBezierCubicCalc']
pub fn im_bezier_cubic_calc(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, t f32)

@[c: 'igImBezierCubicClosestPoint']
pub fn im_bezier_cubic_closest_point(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, p ImVec2, num_segments int)

@[c: 'igImBezierCubicClosestPointCasteljau']
pub fn im_bezier_cubic_closest_point_casteljau(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, p4 ImVec2, p ImVec2, tess_tol f32)

@[c: 'igImBezierQuadraticCalc']
pub fn im_bezier_quadratic_calc(p_out &ImVec2, p1 ImVec2, p2 ImVec2, p3 ImVec2, t f32)

@[c: 'igImLineClosestPoint']
pub fn im_line_closest_point(p_out &ImVec2, a ImVec2, b ImVec2, p ImVec2)

@[c: 'igImTriangleContainsPoint']
pub fn im_triangle_contains_point(a ImVec2, b ImVec2, c ImVec2, p ImVec2) bool

@[c: 'igImTriangleClosestPoint']
pub fn im_triangle_closest_point(p_out &ImVec2, a ImVec2, b ImVec2, c ImVec2, p ImVec2)

@[c: 'igImTriangleBarycentricCoords']
pub fn im_triangle_barycentric_coords(a ImVec2, b ImVec2, c ImVec2, p ImVec2, out_u &f32, out_v &f32, out_w &f32)

@[c: 'igImTriangleArea']
pub fn im_triangle_area(a ImVec2, b ImVec2, c ImVec2) f32

@[c: 'igImTriangleIsClockwise']
pub fn im_triangle_is_clockwise(a ImVec2, b ImVec2, c ImVec2) bool

@[c: 'ImVec1_ImVec1_Nil']
pub fn im_vec1_im_vec1_nil() &ImVec1

@[c: 'ImVec1_destroy']
pub fn im_vec1_destroy(self &ImVec1)

@[c: 'ImVec1_ImVec1_Float']
pub fn im_vec1_im_vec1_float(_x f32) &ImVec1

@[c: 'ImVec2ih_ImVec2ih_Nil']
pub fn im_vec2ih_im_vec2ih_nil() &ImVec2ih

@[c: 'ImVec2ih_destroy']
pub fn im_vec2ih_destroy(self &ImVec2ih)

@[c: 'ImVec2ih_ImVec2ih_short']
pub fn im_vec2ih_im_vec2ih_short(_x i16, _y i16) &ImVec2ih

@[c: 'ImVec2ih_ImVec2ih_Vec2']
pub fn im_vec2ih_im_vec2ih_vec2(rhs ImVec2) &ImVec2ih

@[c: 'ImRect_ImRect_Nil']
pub fn im_rect_im_rect_nil() &ImRect

@[c: 'ImRect_destroy']
pub fn im_rect_destroy(self &ImRect)

@[c: 'ImRect_ImRect_Vec2']
pub fn im_rect_im_rect_vec2(min ImVec2, max ImVec2) &ImRect

@[c: 'ImRect_ImRect_Vec4']
pub fn im_rect_im_rect_vec4(v ImVec4) &ImRect

@[c: 'ImRect_ImRect_Float']
pub fn im_rect_im_rect_float(x1 f32, y1 f32, x2 f32, y2 f32) &ImRect

@[c: 'ImRect_GetCenter']
pub fn im_rect_get_center(p_out &ImVec2, self &ImRect)

@[c: 'ImRect_GetSize']
pub fn im_rect_get_size(p_out &ImVec2, self &ImRect)

@[c: 'ImRect_GetWidth']
pub fn im_rect_get_width(self &ImRect) f32

@[c: 'ImRect_GetHeight']
pub fn im_rect_get_height(self &ImRect) f32

@[c: 'ImRect_GetArea']
pub fn im_rect_get_area(self &ImRect) f32

@[c: 'ImRect_GetTL']
pub fn im_rect_get_tl(p_out &ImVec2, self &ImRect)

@[c: 'ImRect_GetTR']
pub fn im_rect_get_tr(p_out &ImVec2, self &ImRect)

@[c: 'ImRect_GetBL']
pub fn im_rect_get_bl(p_out &ImVec2, self &ImRect)

@[c: 'ImRect_GetBR']
pub fn im_rect_get_br(p_out &ImVec2, self &ImRect)

@[c: 'ImRect_Contains_Vec2']
pub fn im_rect_contains_vec2(self &ImRect, p ImVec2) bool

@[c: 'ImRect_Contains_Rect']
pub fn im_rect_contains_rect(self &ImRect, r ImRect) bool

@[c: 'ImRect_ContainsWithPad']
pub fn im_rect_contains_with_pad(self &ImRect, p ImVec2, pad ImVec2) bool

@[c: 'ImRect_Overlaps']
pub fn im_rect_overlaps(self &ImRect, r ImRect) bool

@[c: 'ImRect_Add_Vec2']
pub fn im_rect_add_vec2(self &ImRect, p ImVec2)

@[c: 'ImRect_Add_Rect']
pub fn im_rect_add_rect(self &ImRect, r ImRect)

@[c: 'ImRect_Expand_Float']
pub fn im_rect_expand_float(self &ImRect, amount f32)

@[c: 'ImRect_Expand_Vec2']
pub fn im_rect_expand_vec2(self &ImRect, amount ImVec2)

@[c: 'ImRect_Translate']
pub fn im_rect_translate(self &ImRect, d ImVec2)

@[c: 'ImRect_TranslateX']
pub fn im_rect_translate_x(self &ImRect, dx f32)

@[c: 'ImRect_TranslateY']
pub fn im_rect_translate_y(self &ImRect, dy f32)

@[c: 'ImRect_ClipWith']
pub fn im_rect_clip_with(self &ImRect, r ImRect)

@[c: 'ImRect_ClipWithFull']
pub fn im_rect_clip_with_full(self &ImRect, r ImRect)

@[c: 'ImRect_Floor']
pub fn im_rect_floor(self &ImRect)

@[c: 'ImRect_IsInverted']
pub fn im_rect_is_inverted(self &ImRect) bool

@[c: 'ImRect_ToVec4']
pub fn im_rect_to_vec4(p_out &ImVec4, self &ImRect)

@[c: 'igImBitArrayGetStorageSizeInBytes']
pub fn im_bit_array_get_storage_size_in_bytes(bitcount int) usize

@[c: 'igImBitArrayClearAllBits']
pub fn im_bit_array_clear_all_bits(arr &ImU32, bitcount int)

@[c: 'igImBitArrayTestBit']
pub fn im_bit_array_test_bit(arr &ImU32, n int) bool

@[c: 'igImBitArrayClearBit']
pub fn im_bit_array_clear_bit(arr &ImU32, n int)

@[c: 'igImBitArraySetBit']
pub fn im_bit_array_set_bit(arr &ImU32, n int)

@[c: 'igImBitArraySetBitRange']
pub fn im_bit_array_set_bit_range(arr &ImU32, n int, n2 int)

@[c: 'ImBitVector_Create']
pub fn im_bit_vector_create(self &ImBitVector, sz int)

@[c: 'ImBitVector_Clear']
pub fn im_bit_vector_clear(self &ImBitVector)

@[c: 'ImBitVector_TestBit']
pub fn im_bit_vector_test_bit(self &ImBitVector, n int) bool

@[c: 'ImBitVector_SetBit']
pub fn im_bit_vector_set_bit(self &ImBitVector, n int)

@[c: 'ImBitVector_ClearBit']
pub fn im_bit_vector_clear_bit(self &ImBitVector, n int)

@[c: 'TextIndex_clear']
pub fn text_index_clear(self &TextIndex)

@[c: 'TextIndex_size']
pub fn text_index_size(self &TextIndex) int

@[c: 'TextIndex_get_line_begin']
pub fn text_index_get_line_begin(self &TextIndex, base &i8, n int) &i8

@[c: 'TextIndex_get_line_end']
pub fn text_index_get_line_end(self &TextIndex, base &i8, n int) &i8

@[c: 'TextIndex_append']
pub fn text_index_append(self &TextIndex, base &i8, old_size int, new_size int)

@[c: 'igImLowerBound']
pub fn im_lower_bound(in_begin &StoragePair, in_end &StoragePair, key ID) &StoragePair

@[c: 'ImDrawListSharedData_ImDrawListSharedData']
pub fn im_draw_list_shared_data_im_draw_list_shared_data() &ImDrawListSharedData

@[c: 'ImDrawListSharedData_destroy']
pub fn im_draw_list_shared_data_destroy(self &ImDrawListSharedData)

@[c: 'ImDrawListSharedData_SetCircleTessellationMaxError']
pub fn im_draw_list_shared_data_set_circle_tessellation_max_error(self &ImDrawListSharedData, max_error f32)

@[c: 'ImDrawDataBuilder_ImDrawDataBuilder']
pub fn im_draw_data_builder_im_draw_data_builder() &ImDrawDataBuilder

@[c: 'ImDrawDataBuilder_destroy']
pub fn im_draw_data_builder_destroy(self &ImDrawDataBuilder)

@[c: 'StyleVarInfo_GetVarPtr']
pub fn style_var_info_get_var_ptr(self &StyleVarInfo, parent voidptr) voidptr

@[c: 'StyleMod_StyleMod_Int']
pub fn style_mod_im_gui_style_mod_int(idx StyleVar, v int) &StyleMod

@[c: 'StyleMod_destroy']
pub fn style_mod_destroy(self &StyleMod)

@[c: 'StyleMod_StyleMod_Float']
pub fn style_mod_im_gui_style_mod_float(idx StyleVar, v f32) &StyleMod

@[c: 'StyleMod_StyleMod_Vec2']
pub fn style_mod_im_gui_style_mod_vec2(idx StyleVar, v ImVec2) &StyleMod

@[c: 'ComboPreviewData_ComboPreviewData']
pub fn combo_preview_data_im_gui_combo_preview_data() &ComboPreviewData

@[c: 'ComboPreviewData_destroy']
pub fn combo_preview_data_destroy(self &ComboPreviewData)

@[c: 'MenuColumns_MenuColumns']
pub fn menu_columns_im_gui_menu_columns() &MenuColumns

@[c: 'MenuColumns_destroy']
pub fn menu_columns_destroy(self &MenuColumns)

@[c: 'MenuColumns_Update']
pub fn menu_columns_update(self &MenuColumns, spacing f32, window_reappearing bool)

@[c: 'MenuColumns_DeclColumns']
pub fn menu_columns_decl_columns(self &MenuColumns, w_icon f32, w_label f32, w_shortcut f32, w_mark f32) f32

@[c: 'MenuColumns_CalcNextTotalWidth']
pub fn menu_columns_calc_next_total_width(self &MenuColumns, update_offsets bool)

@[c: 'InputTextDeactivatedState_InputTextDeactivatedState']
pub fn input_text_deactivated_state_im_gui_input_text_deactivated_state() &InputTextDeactivatedState

@[c: 'InputTextDeactivatedState_destroy']
pub fn input_text_deactivated_state_destroy(self &InputTextDeactivatedState)

@[c: 'InputTextDeactivatedState_ClearFreeMemory']
pub fn input_text_deactivated_state_clear_free_memory(self &InputTextDeactivatedState)

@[c: 'InputTextState_InputTextState']
pub fn input_text_state_im_gui_input_text_state() &InputTextState

@[c: 'InputTextState_destroy']
pub fn input_text_state_destroy(self &InputTextState)

@[c: 'InputTextState_ClearText']
pub fn input_text_state_clear_text(self &InputTextState)

@[c: 'InputTextState_ClearFreeMemory']
pub fn input_text_state_clear_free_memory(self &InputTextState)

@[c: 'InputTextState_OnKeyPressed']
pub fn input_text_state_on_key_pressed(self &InputTextState, key int)

@[c: 'InputTextState_OnCharPressed']
pub fn input_text_state_on_char_pressed(self &InputTextState, c u32)

@[c: 'InputTextState_CursorAnimReset']
pub fn input_text_state_cursor_anim_reset(self &InputTextState)

@[c: 'InputTextState_CursorClamp']
pub fn input_text_state_cursor_clamp(self &InputTextState)

@[c: 'InputTextState_HasSelection']
pub fn input_text_state_has_selection(self &InputTextState) bool

@[c: 'InputTextState_ClearSelection']
pub fn input_text_state_clear_selection(self &InputTextState)

@[c: 'InputTextState_GetCursorPos']
pub fn input_text_state_get_cursor_pos(self &InputTextState) int

@[c: 'InputTextState_GetSelectionStart']
pub fn input_text_state_get_selection_start(self &InputTextState) int

@[c: 'InputTextState_GetSelectionEnd']
pub fn input_text_state_get_selection_end(self &InputTextState) int

@[c: 'InputTextState_SelectAll']
pub fn input_text_state_select_all(self &InputTextState)

@[c: 'InputTextState_ReloadUserBufAndSelectAll']
pub fn input_text_state_reload_user_buf_and_select_all(self &InputTextState)

@[c: 'InputTextState_ReloadUserBufAndKeepSelection']
pub fn input_text_state_reload_user_buf_and_keep_selection(self &InputTextState)

@[c: 'InputTextState_ReloadUserBufAndMoveToEnd']
pub fn input_text_state_reload_user_buf_and_move_to_end(self &InputTextState)

@[c: 'NextWindowData_NextWindowData']
pub fn next_window_data_im_gui_next_window_data() &NextWindowData

@[c: 'NextWindowData_destroy']
pub fn next_window_data_destroy(self &NextWindowData)

@[c: 'NextWindowData_ClearFlags']
pub fn next_window_data_clear_flags(self &NextWindowData)

@[c: 'NextItemData_NextItemData']
pub fn next_item_data_im_gui_next_item_data() &NextItemData

@[c: 'NextItemData_destroy']
pub fn next_item_data_destroy(self &NextItemData)

@[c: 'NextItemData_ClearFlags']
pub fn next_item_data_clear_flags(self &NextItemData)

@[c: 'LastItemData_LastItemData']
pub fn last_item_data_im_gui_last_item_data() &LastItemData

@[c: 'LastItemData_destroy']
pub fn last_item_data_destroy(self &LastItemData)

@[c: 'ErrorRecoveryState_ErrorRecoveryState']
pub fn error_recovery_state_im_gui_error_recovery_state() &ErrorRecoveryState

@[c: 'ErrorRecoveryState_destroy']
pub fn error_recovery_state_destroy(self &ErrorRecoveryState)

@[c: 'PtrOrIndex_PtrOrIndex_Ptr']
pub fn ptr_or_index_im_gui_ptr_or_index_ptr(ptr voidptr) &PtrOrIndex

@[c: 'PtrOrIndex_destroy']
pub fn ptr_or_index_destroy(self &PtrOrIndex)

@[c: 'PtrOrIndex_PtrOrIndex_Int']
pub fn ptr_or_index_im_gui_ptr_or_index_int(index int) &PtrOrIndex

@[c: 'PopupData_PopupData']
pub fn popup_data_im_gui_popup_data() &PopupData

@[c: 'PopupData_destroy']
pub fn popup_data_destroy(self &PopupData)

@[c: 'InputEvent_InputEvent']
pub fn input_event_im_gui_input_event() &InputEvent

@[c: 'InputEvent_destroy']
pub fn input_event_destroy(self &InputEvent)

@[c: 'KeyRoutingData_KeyRoutingData']
pub fn key_routing_data_im_gui_key_routing_data() &KeyRoutingData

@[c: 'KeyRoutingData_destroy']
pub fn key_routing_data_destroy(self &KeyRoutingData)

@[c: 'KeyRoutingTable_KeyRoutingTable']
pub fn key_routing_table_im_gui_key_routing_table() &KeyRoutingTable

@[c: 'KeyRoutingTable_destroy']
pub fn key_routing_table_destroy(self &KeyRoutingTable)

@[c: 'KeyRoutingTable_Clear']
pub fn key_routing_table_clear(self &KeyRoutingTable)

@[c: 'KeyOwnerData_KeyOwnerData']
pub fn key_owner_data_im_gui_key_owner_data() &KeyOwnerData

@[c: 'KeyOwnerData_destroy']
pub fn key_owner_data_destroy(self &KeyOwnerData)

@[c: 'ListClipperRange_FromIndices']
pub fn list_clipper_range_from_indices(min int, max int) ListClipperRange

@[c: 'ListClipperRange_FromPositions']
pub fn list_clipper_range_from_positions(y1 f32, y2 f32, off_min int, off_max int) ListClipperRange

@[c: 'ListClipperData_ListClipperData']
pub fn list_clipper_data_im_gui_list_clipper_data() &ListClipperData

@[c: 'ListClipperData_destroy']
pub fn list_clipper_data_destroy(self &ListClipperData)

@[c: 'ListClipperData_Reset']
pub fn list_clipper_data_reset(self &ListClipperData, clipper &ListClipper)

@[c: 'NavItemData_NavItemData']
pub fn nav_item_data_im_gui_nav_item_data() &NavItemData

@[c: 'NavItemData_destroy']
pub fn nav_item_data_destroy(self &NavItemData)

@[c: 'NavItemData_Clear']
pub fn nav_item_data_clear(self &NavItemData)

@[c: 'TypingSelectState_TypingSelectState']
pub fn typing_select_state_im_gui_typing_select_state() &TypingSelectState

@[c: 'TypingSelectState_destroy']
pub fn typing_select_state_destroy(self &TypingSelectState)

@[c: 'TypingSelectState_Clear']
pub fn typing_select_state_clear(self &TypingSelectState)

@[c: 'OldColumnData_OldColumnData']
pub fn old_column_data_im_gui_old_column_data() &OldColumnData

@[c: 'OldColumnData_destroy']
pub fn old_column_data_destroy(self &OldColumnData)

@[c: 'OldColumns_OldColumns']
pub fn old_columns_im_gui_old_columns() &OldColumns

@[c: 'OldColumns_destroy']
pub fn old_columns_destroy(self &OldColumns)

@[c: 'BoxSelectState_BoxSelectState']
pub fn box_select_state_im_gui_box_select_state() &BoxSelectState

@[c: 'BoxSelectState_destroy']
pub fn box_select_state_destroy(self &BoxSelectState)

@[c: 'MultiSelectTempData_MultiSelectTempData']
pub fn multi_select_temp_data_im_gui_multi_select_temp_data() &MultiSelectTempData

@[c: 'MultiSelectTempData_destroy']
pub fn multi_select_temp_data_destroy(self &MultiSelectTempData)

@[c: 'MultiSelectTempData_Clear']
pub fn multi_select_temp_data_clear(self &MultiSelectTempData)

@[c: 'MultiSelectTempData_ClearIO']
pub fn multi_select_temp_data_clear_io(self &MultiSelectTempData)

@[c: 'MultiSelectState_MultiSelectState']
pub fn multi_select_state_im_gui_multi_select_state() &MultiSelectState

@[c: 'MultiSelectState_destroy']
pub fn multi_select_state_destroy(self &MultiSelectState)

@[c: 'DockNode_DockNode']
pub fn dock_node_im_gui_dock_node(id ID) &DockNode

@[c: 'DockNode_destroy']
pub fn dock_node_destroy(self &DockNode)

@[c: 'DockNode_IsRootNode']
pub fn dock_node_is_root_node(self &DockNode) bool

@[c: 'DockNode_IsDockSpace']
pub fn dock_node_is_dock_space(self &DockNode) bool

@[c: 'DockNode_IsFloatingNode']
pub fn dock_node_is_floating_node(self &DockNode) bool

@[c: 'DockNode_IsCentralNode']
pub fn dock_node_is_central_node(self &DockNode) bool

@[c: 'DockNode_IsHiddenTabBar']
pub fn dock_node_is_hidden_tab_bar(self &DockNode) bool

@[c: 'DockNode_IsNoTabBar']
pub fn dock_node_is_no_tab_bar(self &DockNode) bool

@[c: 'DockNode_IsSplitNode']
pub fn dock_node_is_split_node(self &DockNode) bool

@[c: 'DockNode_IsLeafNode']
pub fn dock_node_is_leaf_node(self &DockNode) bool

@[c: 'DockNode_IsEmpty']
pub fn dock_node_is_empty(self &DockNode) bool

@[c: 'DockNode_Rect']
pub fn dock_node_rect(p_out &ImRect, self &DockNode)

@[c: 'DockNode_SetLocalFlags']
pub fn dock_node_set_local_flags(self &DockNode, flags DockNodeFlags)

@[c: 'DockNode_UpdateMergedFlags']
pub fn dock_node_update_merged_flags(self &DockNode)

@[c: 'DockContext_DockContext']
pub fn dock_context_im_gui_dock_context() &DockContext

@[c: 'DockContext_destroy']
pub fn dock_context_destroy(self &DockContext)

@[c: 'ViewportP_ViewportP']
pub fn viewport_p_im_gui_viewport_p() &ViewportP

@[c: 'ViewportP_destroy']
pub fn viewport_p_destroy(self &ViewportP)

@[c: 'ViewportP_ClearRequestFlags']
pub fn viewport_p_clear_request_flags(self &ViewportP)

@[c: 'ViewportP_CalcWorkRectPos']
pub fn viewport_p_calc_work_rect_pos(p_out &ImVec2, self &ViewportP, inset_min ImVec2)

@[c: 'ViewportP_CalcWorkRectSize']
pub fn viewport_p_calc_work_rect_size(p_out &ImVec2, self &ViewportP, inset_min ImVec2, inset_max ImVec2)

@[c: 'ViewportP_UpdateWorkRect']
pub fn viewport_p_update_work_rect(self &ViewportP)

@[c: 'ViewportP_GetMainRect']
pub fn viewport_p_get_main_rect(p_out &ImRect, self &ViewportP)

@[c: 'ViewportP_GetWorkRect']
pub fn viewport_p_get_work_rect(p_out &ImRect, self &ViewportP)

@[c: 'ViewportP_GetBuildWorkRect']
pub fn viewport_p_get_build_work_rect(p_out &ImRect, self &ViewportP)

@[c: 'WindowSettings_WindowSettings']
pub fn window_settings_im_gui_window_settings() &WindowSettings

@[c: 'WindowSettings_destroy']
pub fn window_settings_destroy(self &WindowSettings)

@[c: 'WindowSettings_GetName']
pub fn window_settings_get_name(self &WindowSettings) &i8

@[c: 'SettingsHandler_SettingsHandler']
pub fn settings_handler_im_gui_settings_handler() &SettingsHandler

@[c: 'SettingsHandler_destroy']
pub fn settings_handler_destroy(self &SettingsHandler)

@[c: 'DebugAllocInfo_DebugAllocInfo']
pub fn debug_alloc_info_im_gui_debug_alloc_info() &DebugAllocInfo

@[c: 'DebugAllocInfo_destroy']
pub fn debug_alloc_info_destroy(self &DebugAllocInfo)

@[c: 'StackLevelInfo_StackLevelInfo']
pub fn stack_level_info_im_gui_stack_level_info() &StackLevelInfo

@[c: 'StackLevelInfo_destroy']
pub fn stack_level_info_destroy(self &StackLevelInfo)

@[c: 'IDStackTool_IDStackTool']
pub fn ids_tack_tool_im_gui_ids_tack_tool() &IDStackTool

@[c: 'IDStackTool_destroy']
pub fn ids_tack_tool_destroy(self &IDStackTool)

@[c: 'ContextHook_ContextHook']
pub fn context_hook_im_gui_context_hook() &ContextHook

@[c: 'ContextHook_destroy']
pub fn context_hook_destroy(self &ContextHook)

@[c: 'Context_Context']
pub fn context_im_gui_context(shared_font_atlas &ImFontAtlas) &Context

@[c: 'Context_destroy']
pub fn context_destroy(self &Context)

@[c: 'Window_Window']
pub fn window_im_gui_window(context &Context, name &i8) &Window

@[c: 'Window_destroy']
pub fn window_destroy(self &Window)

@[c: 'Window_GetID_Str']
pub fn window_get_id_str(self &Window, str &i8, str_end &i8) ID

@[c: 'Window_GetID_Ptr']
pub fn window_get_id_ptr(self &Window, ptr voidptr) ID

@[c: 'Window_GetID_Int']
pub fn window_get_id_int(self &Window, n int) ID

@[c: 'Window_GetIDFromPos']
pub fn window_get_idf_rom_pos(self &Window, p_abs ImVec2) ID

@[c: 'Window_GetIDFromRectangle']
pub fn window_get_idf_rom_rectangle(self &Window, r_abs ImRect) ID

@[c: 'Window_Rect']
pub fn window_rect(p_out &ImRect, self &Window)

@[c: 'Window_CalcFontSize']
pub fn window_calc_font_size(self &Window) f32

@[c: 'Window_TitleBarRect']
pub fn window_title_bar_rect(p_out &ImRect, self &Window)

@[c: 'Window_MenuBarRect']
pub fn window_menu_bar_rect(p_out &ImRect, self &Window)

@[c: 'TabItem_TabItem']
pub fn tab_item_im_gui_tab_item() &TabItem

@[c: 'TabItem_destroy']
pub fn tab_item_destroy(self &TabItem)

@[c: 'TabBar_TabBar']
pub fn tab_bar_im_gui_tab_bar() &TabBar

@[c: 'TabBar_destroy']
pub fn tab_bar_destroy(self &TabBar)

@[c: 'TableColumn_TableColumn']
pub fn table_column_im_gui_table_column() &TableColumn

@[c: 'TableColumn_destroy']
pub fn table_column_destroy(self &TableColumn)

@[c: 'TableInstanceData_TableInstanceData']
pub fn table_instance_data_im_gui_table_instance_data() &TableInstanceData

@[c: 'TableInstanceData_destroy']
pub fn table_instance_data_destroy(self &TableInstanceData)

@[c: 'Table_Table']
pub fn table_im_gui_table() &Table

@[c: 'Table_destroy']
pub fn table_destroy(self &Table)

@[c: 'TableTempData_TableTempData']
pub fn table_temp_data_im_gui_table_temp_data() &TableTempData

@[c: 'TableTempData_destroy']
pub fn table_temp_data_destroy(self &TableTempData)

@[c: 'TableColumnSettings_TableColumnSettings']
pub fn table_column_settings_im_gui_table_column_settings() &TableColumnSettings

@[c: 'TableColumnSettings_destroy']
pub fn table_column_settings_destroy(self &TableColumnSettings)

@[c: 'TableSettings_TableSettings']
pub fn table_settings_im_gui_table_settings() &TableSettings

@[c: 'TableSettings_destroy']
pub fn table_settings_destroy(self &TableSettings)

@[c: 'TableSettings_GetColumnSettings']
pub fn table_settings_get_column_settings(self &TableSettings) &TableColumnSettings

@[c: 'igGetIO_ContextPtr']
pub fn get_io_context_ptr(ctx &Context) &IO

@[c: 'igGetPlatformIO_ContextPtr']
pub fn get_platform_io_context_ptr(ctx &Context) &PlatformIO

@[c: 'igGetCurrentWindowRead']
pub fn get_current_window_read() &Window

@[c: 'igGetCurrentWindow']
pub fn get_current_window() &Window

@[c: 'igFindWindowByID']
pub fn find_window_by_id(id ID) &Window

@[c: 'igFindWindowByName']
pub fn find_window_by_name(name &i8) &Window

@[c: 'igUpdateWindowParentAndRootLinks']
pub fn update_window_parent_and_root_links(window &Window, flags WindowFlags, parent_window &Window)

@[c: 'igUpdateWindowSkipRefresh']
pub fn update_window_skip_refresh(window &Window)

@[c: 'igCalcWindowNextAutoFitSize']
pub fn calc_window_next_auto_fit_size(p_out &ImVec2, window &Window)

@[c: 'igIsWindowChildOf']
pub fn is_window_child_of(window &Window, potential_parent &Window, popup_hierarchy bool, dock_hierarchy bool) bool

@[c: 'igIsWindowWithinBeginStackOf']
pub fn is_window_within_begin_stack_of(window &Window, potential_parent &Window) bool

@[c: 'igIsWindowAbove']
pub fn is_window_above(potential_above &Window, potential_below &Window) bool

@[c: 'igIsWindowNavFocusable']
pub fn is_window_nav_focusable(window &Window) bool

@[c: 'igSetWindowPos_WindowPtr']
pub fn set_window_pos_window_ptr(window &Window, pos ImVec2, cond Cond)

@[c: 'igSetWindowSize_WindowPtr']
pub fn set_window_size_window_ptr(window &Window, size ImVec2, cond Cond)

@[c: 'igSetWindowCollapsed_WindowPtr']
pub fn set_window_collapsed_window_ptr(window &Window, collapsed bool, cond Cond)

@[c: 'igSetWindowHitTestHole']
pub fn set_window_hit_test_hole(window &Window, pos ImVec2, size ImVec2)

@[c: 'igSetWindowHiddenAndSkipItemsForCurrentFrame']
pub fn set_window_hidden_and_skip_items_for_current_frame(window &Window)

@[c: 'igSetWindowParentWindowForFocusRoute']
pub fn set_window_parent_window_for_focus_route(window &Window, parent_window &Window)

@[c: 'igWindowRectAbsToRel']
pub fn window_rect_abs_to_rel(p_out &ImRect, window &Window, r ImRect)

@[c: 'igWindowRectRelToAbs']
pub fn window_rect_rel_to_abs(p_out &ImRect, window &Window, r ImRect)

@[c: 'igWindowPosAbsToRel']
pub fn window_pos_abs_to_rel(p_out &ImVec2, window &Window, p ImVec2)

@[c: 'igWindowPosRelToAbs']
pub fn window_pos_rel_to_abs(p_out &ImVec2, window &Window, p ImVec2)

@[c: 'igFocusWindow']
pub fn focus_window(window &Window, flags FocusRequestFlags)

@[c: 'igFocusTopMostWindowUnderOne']
pub fn focus_top_most_window_under_one(under_this_window &Window, ignore_window &Window, filter_viewport &Viewport, flags FocusRequestFlags)

@[c: 'igBringWindowToFocusFront']
pub fn bring_window_to_focus_front(window &Window)

@[c: 'igBringWindowToDisplayFront']
pub fn bring_window_to_display_front(window &Window)

@[c: 'igBringWindowToDisplayBack']
pub fn bring_window_to_display_back(window &Window)

@[c: 'igBringWindowToDisplayBehind']
pub fn bring_window_to_display_behind(window &Window, above_window &Window)

@[c: 'igFindWindowDisplayIndex']
pub fn find_window_display_index(window &Window) int

@[c: 'igFindBottomMostVisibleWindowWithinBeginStack']
pub fn find_bottom_most_visible_window_within_begin_stack(window &Window) &Window

@[c: 'igSetNextWindowRefreshPolicy']
pub fn set_next_window_refresh_policy(flags WindowRefreshFlags)

@[c: 'igSetCurrentFont']
pub fn set_current_font(font &ImFont)

@[c: 'igGetDefaultFont']
pub fn get_default_font() &ImFont

@[c: 'igPushPasswordFont']
pub fn push_password_font()

@[c: 'igGetForegroundDrawList_WindowPtr']
pub fn get_foreground_draw_list_window_ptr(window &Window) &ImDrawList

@[c: 'igAddDrawListToDrawDataEx']
pub fn add_draw_list_to_draw_data_ex(draw_data &ImDrawData, out_list &ImVector_ImDrawListPtr, draw_list &ImDrawList)

@[c: 'igInitialize']
pub fn initialize()

@[c: 'igShutdown']
pub fn shutdown()

@[c: 'igUpdateInputEvents']
pub fn update_input_events(trickle_fast_inputs bool)

@[c: 'igUpdateHoveredWindowAndCaptureFlags']
pub fn update_hovered_window_and_capture_flags()

@[c: 'igFindHoveredWindowEx']
pub fn find_hovered_window_ex(pos ImVec2, find_first_and_in_any_viewport bool, out_hovered_window &&Window, out_hovered_window_under_moving_window &&Window)

@[c: 'igStartMouseMovingWindow']
pub fn start_mouse_moving_window(window &Window)

@[c: 'igStartMouseMovingWindowOrNode']
pub fn start_mouse_moving_window_or_node(window &Window, node &DockNode, undock bool)

@[c: 'igUpdateMouseMovingWindowNewFrame']
pub fn update_mouse_moving_window_new_frame()

@[c: 'igUpdateMouseMovingWindowEndFrame']
pub fn update_mouse_moving_window_end_frame()

@[c: 'igAddContextHook']
pub fn add_context_hook(context &Context, hook &ContextHook) ID

@[c: 'igRemoveContextHook']
pub fn remove_context_hook(context &Context, hook_to_remove ID)

@[c: 'igCallContextHooks']
pub fn call_context_hooks(context &Context, type_ ContextHookType)

@[c: 'igTranslateWindowsInViewport']
pub fn translate_windows_in_viewport(viewport &ViewportP, old_pos ImVec2, new_pos ImVec2, old_size ImVec2, new_size ImVec2)

@[c: 'igScaleWindowsInViewport']
pub fn scale_windows_in_viewport(viewport &ViewportP, scale f32)

@[c: 'igDestroyPlatformWindow']
pub fn destroy_platform_window(viewport &ViewportP)

@[c: 'igSetWindowViewport']
pub fn set_window_viewport(window &Window, viewport &ViewportP)

@[c: 'igSetCurrentViewport']
pub fn set_current_viewport(window &Window, viewport &ViewportP)

@[c: 'igGetViewportPlatformMonitor']
pub fn get_viewport_platform_monitor(viewport &Viewport) &PlatformMonitor

@[c: 'igFindHoveredViewportFromPlatformWindowStack']
pub fn find_hovered_viewport_from_platform_window_stack(mouse_platform_pos ImVec2) &ViewportP

@[c: 'igMarkIniSettingsDirty_Nil']
pub fn mark_ini_settings_dirty_nil()

@[c: 'igMarkIniSettingsDirty_WindowPtr']
pub fn mark_ini_settings_dirty_window_ptr(window &Window)

@[c: 'igClearIniSettings']
pub fn clear_ini_settings()

@[c: 'igAddSettingsHandler']
pub fn add_settings_handler(handler &SettingsHandler)

@[c: 'igRemoveSettingsHandler']
pub fn remove_settings_handler(type_name &i8)

@[c: 'igFindSettingsHandler']
pub fn find_settings_handler(type_name &i8) &SettingsHandler

@[c: 'igCreateNewWindowSettings']
pub fn create_new_window_settings(name &i8) &WindowSettings

@[c: 'igFindWindowSettingsByID']
pub fn find_window_settings_by_id(id ID) &WindowSettings

@[c: 'igFindWindowSettingsByWindow']
pub fn find_window_settings_by_window(window &Window) &WindowSettings

@[c: 'igClearWindowSettings']
pub fn clear_window_settings(name &i8)

@[c: 'igLocalizeRegisterEntries']
pub fn localize_register_entries(entries &LocEntry, count int)

@[c: 'igLocalizeGetMsg']
pub fn localize_get_msg(key LocKey) &i8

@[c: 'igSetScrollX_WindowPtr']
pub fn set_scroll_x_window_ptr(window &Window, scroll_x f32)

@[c: 'igSetScrollY_WindowPtr']
pub fn set_scroll_y_window_ptr(window &Window, scroll_y f32)

@[c: 'igSetScrollFromPosX_WindowPtr']
pub fn set_scroll_from_pos_x_window_ptr(window &Window, local_x f32, center_x_ratio f32)

@[c: 'igSetScrollFromPosY_WindowPtr']
pub fn set_scroll_from_pos_y_window_ptr(window &Window, local_y f32, center_y_ratio f32)

@[c: 'igScrollToItem']
pub fn scroll_to_item(flags ScrollFlags)

@[c: 'igScrollToRect']
pub fn scroll_to_rect(window &Window, rect ImRect, flags ScrollFlags)

@[c: 'igScrollToRectEx']
pub fn scroll_to_rect_ex(p_out &ImVec2, window &Window, rect ImRect, flags ScrollFlags)

@[c: 'igScrollToBringRectIntoView']
pub fn scroll_to_bring_rect_into_view(window &Window, rect ImRect)

@[c: 'igGetItemStatusFlags']
pub fn get_item_status_flags() ItemStatusFlags

@[c: 'igGetItemFlags']
pub fn get_item_flags() ItemFlags

@[c: 'igGetActiveID']
pub fn get_active_id() ID

@[c: 'igGetFocusID']
pub fn get_focus_id() ID

@[c: 'igSetActiveID']
pub fn set_active_id(id ID, window &Window)

@[c: 'igSetFocusID']
pub fn set_focus_id(id ID, window &Window)

@[c: 'igClearActiveID']
pub fn clear_active_id()

@[c: 'igGetHoveredID']
pub fn get_hovered_id() ID

@[c: 'igSetHoveredID']
pub fn set_hovered_id(id ID)

@[c: 'igKeepAliveID']
pub fn keep_alive_id(id ID)

@[c: 'igMarkItemEdited']
pub fn mark_item_edited(id ID)

@[c: 'igPushOverrideID']
pub fn push_override_id(id ID)

@[c: 'igGetIDWithSeed_Str']
pub fn get_idw_ith_seed_str(str_id_begin &i8, str_id_end &i8, seed ID) ID

@[c: 'igGetIDWithSeed_Int']
pub fn get_idw_ith_seed_int(n int, seed ID) ID

@[c: 'igItemSize_Vec2']
pub fn item_size_vec2(size ImVec2, text_baseline_y f32)

@[c: 'igItemSize_Rect']
pub fn item_size_rect(bb ImRect, text_baseline_y f32)

@[c: 'igItemAdd']
pub fn item_add(bb ImRect, id ID, nav_bb &ImRect, extra_flags ItemFlags) bool

@[c: 'igItemHoverable']
pub fn item_hoverable(bb ImRect, id ID, item_flags ItemFlags) bool

@[c: 'igIsWindowContentHoverable']
pub fn is_window_content_hoverable(window &Window, flags HoveredFlags) bool

@[c: 'igIsClippedEx']
pub fn is_clipped_ex(bb ImRect, id ID) bool

@[c: 'igSetLastItemData']
pub fn set_last_item_data(item_id ID, item_flags ItemFlags, status_flags ItemStatusFlags, item_rect ImRect)

@[c: 'igCalcItemSize']
pub fn calc_item_size(p_out &ImVec2, size ImVec2, default_w f32, default_h f32)

@[c: 'igCalcWrapWidthForPos']
pub fn calc_wrap_width_for_pos(pos ImVec2, wrap_pos_x f32) f32

@[c: 'igPushMultiItemsWidths']
pub fn push_multi_items_widths(components int, width_full f32)

@[c: 'igShrinkWidths']
pub fn shrink_widths(items &ShrinkWidthItem, count int, width_excess f32)

@[c: 'igGetStyleVarInfo']
pub fn get_style_var_info(idx StyleVar) &StyleVarInfo

@[c: 'igBeginDisabledOverrideReenable']
pub fn begin_disabled_override_reenable()

@[c: 'igEndDisabledOverrideReenable']
pub fn end_disabled_override_reenable()

@[c: 'igLogBegin']
pub fn log_begin(flags LogFlags, auto_open_depth int)

@[c: 'igLogToBuffer']
pub fn log_to_buffer(auto_open_depth int)

@[c: 'igLogRenderedText']
pub fn log_rendered_text(ref_pos &ImVec2, text &i8, text_end &i8)

@[c: 'igLogSetNextTextDecoration']
pub fn log_set_next_text_decoration(prefix &i8, suffix &i8)

@[c: 'igBeginChildEx']
pub fn begin_child_ex(name &i8, id ID, size_arg ImVec2, child_flags ChildFlags, window_flags WindowFlags) bool

@[c: 'igBeginPopupEx']
pub fn begin_popup_ex(id ID, extra_window_flags WindowFlags) bool

@[c: 'igBeginPopupMenuEx']
pub fn begin_popup_menu_ex(id ID, label &i8, extra_window_flags WindowFlags) bool

@[c: 'igOpenPopupEx']
pub fn open_popup_ex(id ID, popup_flags PopupFlags)

@[c: 'igClosePopupToLevel']
pub fn close_popup_to_level(remaining int, restore_focus_to_window_under_popup bool)

@[c: 'igClosePopupsOverWindow']
pub fn close_popups_over_window(ref_window &Window, restore_focus_to_window_under_popup bool)

@[c: 'igClosePopupsExceptModals']
pub fn close_popups_except_modals()

@[c: 'igIsPopupOpen_ID']
pub fn is_popup_open_id(id ID, popup_flags PopupFlags) bool

@[c: 'igGetPopupAllowedExtentRect']
pub fn get_popup_allowed_extent_rect(p_out &ImRect, window &Window)

@[c: 'igGetTopMostPopupModal']
pub fn get_top_most_popup_modal() &Window

@[c: 'igGetTopMostAndVisiblePopupModal']
pub fn get_top_most_and_visible_popup_modal() &Window

@[c: 'igFindBlockingModal']
pub fn find_blocking_modal(window &Window) &Window

@[c: 'igFindBestWindowPosForPopup']
pub fn find_best_window_pos_for_popup(p_out &ImVec2, window &Window)

@[c: 'igFindBestWindowPosForPopupEx']
pub fn find_best_window_pos_for_popup_ex(p_out &ImVec2, ref_pos ImVec2, size ImVec2, last_dir &Dir, r_outer ImRect, r_avoid ImRect, policy PopupPositionPolicy)

@[c: 'igBeginTooltipEx']
pub fn begin_tooltip_ex(tooltip_flags TooltipFlags, extra_window_flags WindowFlags) bool

@[c: 'igBeginTooltipHidden']
pub fn begin_tooltip_hidden() bool

@[c: 'igBeginViewportSideBar']
pub fn begin_viewport_side_bar(name &i8, viewport &Viewport, dir Dir, size f32, window_flags WindowFlags) bool

@[c: 'igBeginMenuEx']
pub fn begin_menu_ex(label &i8, icon &i8, enabled bool) bool

@[c: 'igMenuItemEx']
pub fn menu_item_ex(label &i8, icon &i8, shortcut &i8, selected bool, enabled bool) bool

@[c: 'igBeginComboPopup']
pub fn begin_combo_popup(popup_id ID, bb ImRect, flags ComboFlags) bool

@[c: 'igBeginComboPreview']
pub fn begin_combo_preview() bool

@[c: 'igEndComboPreview']
pub fn end_combo_preview()

@[c: 'igNavInitWindow']
pub fn nav_init_window(window &Window, force_reinit bool)

@[c: 'igNavInitRequestApplyResult']
pub fn nav_init_request_apply_result()

@[c: 'igNavMoveRequestButNoResultYet']
pub fn nav_move_request_but_no_result_yet() bool

@[c: 'igNavMoveRequestSubmit']
pub fn nav_move_request_submit(move_dir Dir, clip_dir Dir, move_flags NavMoveFlags, scroll_flags ScrollFlags)

@[c: 'igNavMoveRequestForward']
pub fn nav_move_request_forward(move_dir Dir, clip_dir Dir, move_flags NavMoveFlags, scroll_flags ScrollFlags)

@[c: 'igNavMoveRequestResolveWithLastItem']
pub fn nav_move_request_resolve_with_last_item(result &NavItemData)

@[c: 'igNavMoveRequestResolveWithPastTreeNode']
pub fn nav_move_request_resolve_with_past_tree_node(result &NavItemData, tree_node_data &TreeNodeStackData)

@[c: 'igNavMoveRequestCancel']
pub fn nav_move_request_cancel()

@[c: 'igNavMoveRequestApplyResult']
pub fn nav_move_request_apply_result()

@[c: 'igNavMoveRequestTryWrapping']
pub fn nav_move_request_try_wrapping(window &Window, move_flags NavMoveFlags)

@[c: 'igNavHighlightActivated']
pub fn nav_highlight_activated(id ID)

@[c: 'igNavClearPreferredPosForAxis']
pub fn nav_clear_preferred_pos_for_axis(axis Axis)

@[c: 'igSetNavCursorVisibleAfterMove']
pub fn set_nav_cursor_visible_after_move()

@[c: 'igNavUpdateCurrentWindowIsScrollPushableX']
pub fn nav_update_current_window_is_scroll_pushable_x()

@[c: 'igSetNavWindow']
pub fn set_nav_window(window &Window)

@[c: 'igSetNavID']
pub fn set_nav_id(id ID, nav_layer NavLayer, focus_scope_id ID, rect_rel ImRect)

@[c: 'igSetNavFocusScope']
pub fn set_nav_focus_scope(focus_scope_id ID)

@[c: 'igFocusItem']
pub fn focus_item()

@[c: 'igActivateItemByID']
pub fn activate_item_by_id(id ID)

@[c: 'igIsNamedKey']
pub fn is_named_key(key Key) bool

@[c: 'igIsNamedKeyOrMod']
pub fn is_named_key_or_mod(key Key) bool

@[c: 'igIsLegacyKey']
pub fn is_legacy_key(key Key) bool

@[c: 'igIsKeyboardKey']
pub fn is_keyboard_key(key Key) bool

@[c: 'igIsGamepadKey']
pub fn is_gamepad_key(key Key) bool

@[c: 'igIsMouseKey']
pub fn is_mouse_key(key Key) bool

@[c: 'igIsAliasKey']
pub fn is_alias_key(key Key) bool

@[c: 'igIsLRModKey']
pub fn is_lrm_od_key(key Key) bool

@[c: 'igFixupKeyChord']
pub fn fixup_key_chord(key_chord KeyChord) KeyChord

@[c: 'igConvertSingleModFlagToKey']
pub fn convert_single_mod_flag_to_key(key Key) Key

@[c: 'igGetKeyData_ContextPtr']
pub fn get_key_data_context_ptr(ctx &Context, key Key) &KeyData

@[c: 'igGetKeyData_Key']
pub fn get_key_data_key(key Key) &KeyData

@[c: 'igGetKeyChordName']
pub fn get_key_chord_name(key_chord KeyChord) &i8

@[c: 'igMouseButtonToKey']
pub fn mouse_button_to_key(button MouseButton) Key

@[c: 'igIsMouseDragPastThreshold']
pub fn is_mouse_drag_past_threshold(button MouseButton, lock_threshold f32) bool

@[c: 'igGetKeyMagnitude2d']
pub fn get_key_magnitude2d(p_out &ImVec2, key_left Key, key_right Key, key_up Key, key_down Key)

@[c: 'igGetNavTweakPressedAmount']
pub fn get_nav_tweak_pressed_amount(axis Axis) f32

@[c: 'igCalcTypematicRepeatAmount']
pub fn calc_typematic_repeat_amount(t0 f32, t1 f32, repeat_delay f32, repeat_rate f32) int

@[c: 'igGetTypematicRepeatRate']
pub fn get_typematic_repeat_rate(flags InputFlags, repeat_delay &f32, repeat_rate &f32)

@[c: 'igTeleportMousePos']
pub fn teleport_mouse_pos(pos ImVec2)

@[c: 'igSetActiveIdUsingAllKeyboardKeys']
pub fn set_active_id_using_all_keyboard_keys()

@[c: 'igIsActiveIdUsingNavDir']
pub fn is_active_id_using_nav_dir(dir Dir) bool

@[c: 'igGetKeyOwner']
pub fn get_key_owner(key Key) ID

@[c: 'igSetKeyOwner']
pub fn set_key_owner(key Key, owner_id ID, flags InputFlags)

@[c: 'igSetKeyOwnersForKeyChord']
pub fn set_key_owners_for_key_chord(key KeyChord, owner_id ID, flags InputFlags)

@[c: 'igSetItemKeyOwner_InputFlags']
pub fn set_item_key_owner_input_flags(key Key, flags InputFlags)

@[c: 'igTestKeyOwner']
pub fn test_key_owner(key Key, owner_id ID) bool

@[c: 'igGetKeyOwnerData']
pub fn get_key_owner_data(ctx &Context, key Key) &KeyOwnerData

@[c: 'igIsKeyDown_ID']
pub fn is_key_down_id(key Key, owner_id ID) bool

@[c: 'igIsKeyPressed_InputFlags']
pub fn is_key_pressed_input_flags(key Key, flags InputFlags, owner_id ID) bool

@[c: 'igIsKeyReleased_ID']
pub fn is_key_released_id(key Key, owner_id ID) bool

@[c: 'igIsKeyChordPressed_InputFlags']
pub fn is_key_chord_pressed_input_flags(key_chord KeyChord, flags InputFlags, owner_id ID) bool

@[c: 'igIsMouseDown_ID']
pub fn is_mouse_down_id(button MouseButton, owner_id ID) bool

@[c: 'igIsMouseClicked_InputFlags']
pub fn is_mouse_clicked_input_flags(button MouseButton, flags InputFlags, owner_id ID) bool

@[c: 'igIsMouseReleased_ID']
pub fn is_mouse_released_id(button MouseButton, owner_id ID) bool

@[c: 'igIsMouseDoubleClicked_ID']
pub fn is_mouse_double_clicked_id(button MouseButton, owner_id ID) bool

@[c: 'igShortcut_ID']
pub fn shortcut_id(key_chord KeyChord, flags InputFlags, owner_id ID) bool

@[c: 'igSetShortcutRouting']
pub fn set_shortcut_routing(key_chord KeyChord, flags InputFlags, owner_id ID) bool

@[c: 'igTestShortcutRouting']
pub fn test_shortcut_routing(key_chord KeyChord, owner_id ID) bool

@[c: 'igGetShortcutRoutingData']
pub fn get_shortcut_routing_data(key_chord KeyChord) &KeyRoutingData

@[c: 'igDockContextInitialize']
pub fn dock_context_initialize(ctx &Context)

@[c: 'igDockContextShutdown']
pub fn dock_context_shutdown(ctx &Context)

@[c: 'igDockContextClearNodes']
pub fn dock_context_clear_nodes(ctx &Context, root_id ID, clear_settings_refs bool)

@[c: 'igDockContextRebuildNodes']
pub fn dock_context_rebuild_nodes(ctx &Context)

@[c: 'igDockContextNewFrameUpdateUndocking']
pub fn dock_context_new_frame_update_undocking(ctx &Context)

@[c: 'igDockContextNewFrameUpdateDocking']
pub fn dock_context_new_frame_update_docking(ctx &Context)

@[c: 'igDockContextEndFrame']
pub fn dock_context_end_frame(ctx &Context)

@[c: 'igDockContextGenNodeID']
pub fn dock_context_gen_node_id(ctx &Context) ID

@[c: 'igDockContextQueueDock']
pub fn dock_context_queue_dock(ctx &Context, target &Window, target_node &DockNode, payload &Window, split_dir Dir, split_ratio f32, split_outer bool)

@[c: 'igDockContextQueueUndockWindow']
pub fn dock_context_queue_undock_window(ctx &Context, window &Window)

@[c: 'igDockContextQueueUndockNode']
pub fn dock_context_queue_undock_node(ctx &Context, node &DockNode)

@[c: 'igDockContextProcessUndockWindow']
pub fn dock_context_process_undock_window(ctx &Context, window &Window, clear_persistent_docking_ref bool)

@[c: 'igDockContextProcessUndockNode']
pub fn dock_context_process_undock_node(ctx &Context, node &DockNode)

@[c: 'igDockContextCalcDropPosForDocking']
pub fn dock_context_calc_drop_pos_for_docking(target &Window, target_node &DockNode, payload_window &Window, payload_node &DockNode, split_dir Dir, split_outer bool, out_pos &ImVec2) bool

@[c: 'igDockContextFindNodeByID']
pub fn dock_context_find_node_by_id(ctx &Context, id ID) &DockNode

@[c: 'igDockNodeWindowMenuHandler_Default']
pub fn dock_node_window_menu_handler_default(ctx &Context, node &DockNode, tab_bar &TabBar)

@[c: 'igDockNodeBeginAmendTabBar']
pub fn dock_node_begin_amend_tab_bar(node &DockNode) bool

@[c: 'igDockNodeEndAmendTabBar']
pub fn dock_node_end_amend_tab_bar()

@[c: 'igDockNodeGetRootNode']
pub fn dock_node_get_root_node(node &DockNode) &DockNode

@[c: 'igDockNodeIsInHierarchyOf']
pub fn dock_node_is_in_hierarchy_of(node &DockNode, parent &DockNode) bool

@[c: 'igDockNodeGetDepth']
pub fn dock_node_get_depth(node &DockNode) int

@[c: 'igDockNodeGetWindowMenuButtonId']
pub fn dock_node_get_window_menu_button_id(node &DockNode) ID

@[c: 'igGetWindowDockNode']
pub fn get_window_dock_node() &DockNode

@[c: 'igGetWindowAlwaysWantOwnTabBar']
pub fn get_window_always_want_own_tab_bar(window &Window) bool

@[c: 'igBeginDocked']
pub fn begin_docked(window &Window, p_open &bool)

@[c: 'igBeginDockableDragDropSource']
pub fn begin_dockable_drag_drop_source(window &Window)

@[c: 'igBeginDockableDragDropTarget']
pub fn begin_dockable_drag_drop_target(window &Window)

@[c: 'igSetWindowDock']
pub fn set_window_dock(window &Window, dock_id ID, cond Cond)

@[c: 'igDockBuilderDockWindow']
pub fn dock_builder_dock_window(window_name &i8, node_id ID)

@[c: 'igDockBuilderGetNode']
pub fn dock_builder_get_node(node_id ID) &DockNode

@[c: 'igDockBuilderGetCentralNode']
pub fn dock_builder_get_central_node(node_id ID) &DockNode

@[c: 'igDockBuilderAddNode']
pub fn dock_builder_add_node(node_id ID, flags DockNodeFlags) ID

@[c: 'igDockBuilderRemoveNode']
pub fn dock_builder_remove_node(node_id ID)

@[c: 'igDockBuilderRemoveNodeDockedWindows']
pub fn dock_builder_remove_node_docked_windows(node_id ID, clear_settings_refs bool)

@[c: 'igDockBuilderRemoveNodeChildNodes']
pub fn dock_builder_remove_node_child_nodes(node_id ID)

@[c: 'igDockBuilderSetNodePos']
pub fn dock_builder_set_node_pos(node_id ID, pos ImVec2)

@[c: 'igDockBuilderSetNodeSize']
pub fn dock_builder_set_node_size(node_id ID, size ImVec2)

@[c: 'igDockBuilderSplitNode']
pub fn dock_builder_split_node(node_id ID, split_dir Dir, size_ratio_for_node_at_dir f32, out_id_at_dir &ID, out_id_at_opposite_dir &ID) ID

@[c: 'igDockBuilderCopyDockSpace']
pub fn dock_builder_copy_dock_space(src_dockspace_id ID, dst_dockspace_id ID, in_window_remap_pairs &ImVector_const_charPtr)

@[c: 'igDockBuilderCopyNode']
pub fn dock_builder_copy_node(src_node_id ID, dst_node_id ID, out_node_remap_pairs &ImVector_ID)

@[c: 'igDockBuilderCopyWindowSettings']
pub fn dock_builder_copy_window_settings(src_name &i8, dst_name &i8)

@[c: 'igDockBuilderFinish']
pub fn dock_builder_finish(node_id ID)

@[c: 'igPushFocusScope']
pub fn push_focus_scope(id ID)

@[c: 'igPopFocusScope']
pub fn pop_focus_scope()

@[c: 'igGetCurrentFocusScope']
pub fn get_current_focus_scope() ID

@[c: 'igIsDragDropActive']
pub fn is_drag_drop_active() bool

@[c: 'igBeginDragDropTargetCustom']
pub fn begin_drag_drop_target_custom(bb ImRect, id ID) bool

@[c: 'igClearDragDrop']
pub fn clear_drag_drop()

@[c: 'igIsDragDropPayloadBeingAccepted']
pub fn is_drag_drop_payload_being_accepted() bool

@[c: 'igRenderDragDropTargetRect']
pub fn render_drag_drop_target_rect(bb ImRect, item_clip_rect ImRect)

@[c: 'igGetTypingSelectRequest']
pub fn get_typing_select_request(flags TypingSelectFlags) &TypingSelectRequest

@[c: 'igTypingSelectFindMatch']
pub fn typing_select_find_match(req &TypingSelectRequest, items_count int, get_item_name_func fn (voidptr, int) &i8, user_data voidptr, nav_item_idx int) int

@[c: 'igTypingSelectFindNextSingleCharMatch']
pub fn typing_select_find_next_single_char_match(req &TypingSelectRequest, items_count int, get_item_name_func fn (voidptr, int) &i8, user_data voidptr, nav_item_idx int) int

@[c: 'igTypingSelectFindBestLeadingMatch']
pub fn typing_select_find_best_leading_match(req &TypingSelectRequest, items_count int, get_item_name_func fn (voidptr, int) &i8, user_data voidptr) int

@[c: 'igBeginBoxSelect']
pub fn begin_box_select(scope_rect ImRect, window &Window, box_select_id ID, ms_flags MultiSelectFlags) bool

@[c: 'igEndBoxSelect']
pub fn end_box_select(scope_rect ImRect, ms_flags MultiSelectFlags)

@[c: 'igMultiSelectItemHeader']
pub fn multi_select_item_header(id ID, p_selected &bool, p_button_flags &ButtonFlags)

@[c: 'igMultiSelectItemFooter']
pub fn multi_select_item_footer(id ID, p_selected &bool, p_pressed &bool)

@[c: 'igMultiSelectAddSetAll']
pub fn multi_select_add_set_all(ms &MultiSelectTempData, selected bool)

@[c: 'igMultiSelectAddSetRange']
pub fn multi_select_add_set_range(ms &MultiSelectTempData, selected bool, range_dir int, first_item SelectionUserData, last_item SelectionUserData)

@[c: 'igGetBoxSelectState']
pub fn get_box_select_state(id ID) &BoxSelectState

@[c: 'igGetMultiSelectState']
pub fn get_multi_select_state(id ID) &MultiSelectState

@[c: 'igSetWindowClipRectBeforeSetChannel']
pub fn set_window_clip_rect_before_set_channel(window &Window, clip_rect ImRect)

@[c: 'igBeginColumns']
pub fn begin_columns(str_id &i8, count int, flags OldColumnFlags)

@[c: 'igEndColumns']
pub fn end_columns()

@[c: 'igPushColumnClipRect']
pub fn push_column_clip_rect(column_index int)

@[c: 'igPushColumnsBackground']
pub fn push_columns_background()

@[c: 'igPopColumnsBackground']
pub fn pop_columns_background()

@[c: 'igGetColumnsID']
pub fn get_columns_id(str_id &i8, count int) ID

@[c: 'igFindOrCreateColumns']
pub fn find_or_create_columns(window &Window, id ID) &OldColumns

@[c: 'igGetColumnOffsetFromNorm']
pub fn get_column_offset_from_norm(columns &OldColumns, offset_norm f32) f32

@[c: 'igGetColumnNormFromOffset']
pub fn get_column_norm_from_offset(columns &OldColumns, offset f32) f32

@[c: 'igTableOpenContextMenu']
pub fn table_open_context_menu(column_n int)

@[c: 'igTableSetColumnWidth']
pub fn table_set_column_width(column_n int, width f32)

@[c: 'igTableSetColumnSortDirection']
pub fn table_set_column_sort_direction(column_n int, sort_direction SortDirection, append_to_sort_specs bool)

@[c: 'igTableGetHoveredRow']
pub fn table_get_hovered_row() int

@[c: 'igTableGetHeaderRowHeight']
pub fn table_get_header_row_height() f32

@[c: 'igTableGetHeaderAngledMaxLabelWidth']
pub fn table_get_header_angled_max_label_width() f32

@[c: 'igTablePushBackgroundChannel']
pub fn table_push_background_channel()

@[c: 'igTablePopBackgroundChannel']
pub fn table_pop_background_channel()

@[c: 'igTableAngledHeadersRowEx']
pub fn table_angled_headers_row_ex(row_id ID, angle f32, max_label_width f32, data &TableHeaderData, data_count int)

@[c: 'igGetCurrentTable']
pub fn get_current_table() &Table

@[c: 'igTableFindByID']
pub fn table_find_by_id(id ID) &Table

@[c: 'igBeginTableEx']
pub fn begin_table_ex(name &i8, id ID, columns_count int, flags TableFlags, outer_size ImVec2, inner_width f32) bool

@[c: 'igTableBeginInitMemory']
pub fn table_begin_init_memory(table &Table, columns_count int)

@[c: 'igTableBeginApplyRequests']
pub fn table_begin_apply_requests(table &Table)

@[c: 'igTableSetupDrawChannels']
pub fn table_setup_draw_channels(table &Table)

@[c: 'igTableUpdateLayout']
pub fn table_update_layout(table &Table)

@[c: 'igTableUpdateBorders']
pub fn table_update_borders(table &Table)

@[c: 'igTableUpdateColumnsWeightFromWidth']
pub fn table_update_columns_weight_from_width(table &Table)

@[c: 'igTableDrawBorders']
pub fn table_draw_borders(table &Table)

@[c: 'igTableDrawDefaultContextMenu']
pub fn table_draw_default_context_menu(table &Table, flags_for_section_to_display TableFlags)

@[c: 'igTableBeginContextMenuPopup']
pub fn table_begin_context_menu_popup(table &Table) bool

@[c: 'igTableMergeDrawChannels']
pub fn table_merge_draw_channels(table &Table)

@[c: 'igTableGetInstanceData']
pub fn table_get_instance_data(table &Table, instance_no int) &TableInstanceData

@[c: 'igTableGetInstanceID']
pub fn table_get_instance_id(table &Table, instance_no int) ID

@[c: 'igTableSortSpecsSanitize']
pub fn table_sort_specs_sanitize(table &Table)

@[c: 'igTableSortSpecsBuild']
pub fn table_sort_specs_build(table &Table)

@[c: 'igTableGetColumnNextSortDirection']
pub fn table_get_column_next_sort_direction(column &TableColumn) SortDirection

@[c: 'igTableFixColumnSortDirection']
pub fn table_fix_column_sort_direction(table &Table, column &TableColumn)

@[c: 'igTableGetColumnWidthAuto']
pub fn table_get_column_width_auto(table &Table, column &TableColumn) f32

@[c: 'igTableBeginRow']
pub fn table_begin_row(table &Table)

@[c: 'igTableEndRow']
pub fn table_end_row(table &Table)

@[c: 'igTableBeginCell']
pub fn table_begin_cell(table &Table, column_n int)

@[c: 'igTableEndCell']
pub fn table_end_cell(table &Table)

@[c: 'igTableGetCellBgRect']
pub fn table_get_cell_bg_rect(p_out &ImRect, table &Table, column_n int)

@[c: 'igTableGetColumnName_TablePtr']
pub fn table_get_column_name_table_ptr(table &Table, column_n int) &i8

@[c: 'igTableGetColumnResizeID']
pub fn table_get_column_resize_id(table &Table, column_n int, instance_no int) ID

@[c: 'igTableCalcMaxColumnWidth']
pub fn table_calc_max_column_width(table &Table, column_n int) f32

@[c: 'igTableSetColumnWidthAutoSingle']
pub fn table_set_column_width_auto_single(table &Table, column_n int)

@[c: 'igTableSetColumnWidthAutoAll']
pub fn table_set_column_width_auto_all(table &Table)

@[c: 'igTableRemove']
pub fn table_remove(table &Table)

@[c: 'igTableGcCompactTransientBuffers_TablePtr']
pub fn table_gc_compact_transient_buffers_table_ptr(table &Table)

@[c: 'igTableGcCompactTransientBuffers_TableTempDataPtr']
pub fn table_gc_compact_transient_buffers_table_temp_data_ptr(table &TableTempData)

@[c: 'igTableGcCompactSettings']
pub fn table_gc_compact_settings()

@[c: 'igTableLoadSettings']
pub fn table_load_settings(table &Table)

@[c: 'igTableSaveSettings']
pub fn table_save_settings(table &Table)

@[c: 'igTableResetSettings']
pub fn table_reset_settings(table &Table)

@[c: 'igTableGetBoundSettings']
pub fn table_get_bound_settings(table &Table) &TableSettings

@[c: 'igTableSettingsAddSettingsHandler']
pub fn table_settings_add_settings_handler()

@[c: 'igTableSettingsCreate']
pub fn table_settings_create(id ID, columns_count int) &TableSettings

@[c: 'igTableSettingsFindByID']
pub fn table_settings_find_by_id(id ID) &TableSettings

@[c: 'igGetCurrentTabBar']
pub fn get_current_tab_bar() &TabBar

@[c: 'igBeginTabBarEx']
pub fn begin_tab_bar_ex(tab_bar &TabBar, bb ImRect, flags TabBarFlags) bool

@[c: 'igTabBarFindTabByID']
pub fn tab_bar_find_tab_by_id(tab_bar &TabBar, tab_id ID) &TabItem

@[c: 'igTabBarFindTabByOrder']
pub fn tab_bar_find_tab_by_order(tab_bar &TabBar, order int) &TabItem

@[c: 'igTabBarFindMostRecentlySelectedTabForActiveWindow']
pub fn tab_bar_find_most_recently_selected_tab_for_active_window(tab_bar &TabBar) &TabItem

@[c: 'igTabBarGetCurrentTab']
pub fn tab_bar_get_current_tab(tab_bar &TabBar) &TabItem

@[c: 'igTabBarGetTabOrder']
pub fn tab_bar_get_tab_order(tab_bar &TabBar, tab &TabItem) int

@[c: 'igTabBarGetTabName']
pub fn tab_bar_get_tab_name(tab_bar &TabBar, tab &TabItem) &i8

@[c: 'igTabBarAddTab']
pub fn tab_bar_add_tab(tab_bar &TabBar, tab_flags TabItemFlags, window &Window)

@[c: 'igTabBarRemoveTab']
pub fn tab_bar_remove_tab(tab_bar &TabBar, tab_id ID)

@[c: 'igTabBarCloseTab']
pub fn tab_bar_close_tab(tab_bar &TabBar, tab &TabItem)

@[c: 'igTabBarQueueFocus_TabItemPtr']
pub fn tab_bar_queue_focus_tab_item_ptr(tab_bar &TabBar, tab &TabItem)

@[c: 'igTabBarQueueFocus_Str']
pub fn tab_bar_queue_focus_str(tab_bar &TabBar, tab_name &i8)

@[c: 'igTabBarQueueReorder']
pub fn tab_bar_queue_reorder(tab_bar &TabBar, tab &TabItem, offset int)

@[c: 'igTabBarQueueReorderFromMousePos']
pub fn tab_bar_queue_reorder_from_mouse_pos(tab_bar &TabBar, tab &TabItem, mouse_pos ImVec2)

@[c: 'igTabBarProcessReorder']
pub fn tab_bar_process_reorder(tab_bar &TabBar) bool

@[c: 'igTabItemEx']
pub fn tab_item_ex(tab_bar &TabBar, label &i8, p_open &bool, flags TabItemFlags, docked_window &Window) bool

@[c: 'igTabItemSpacing']
pub fn tab_item_spacing(str_id &i8, flags TabItemFlags, width f32)

@[c: 'igTabItemCalcSize_Str']
pub fn tab_item_calc_size_str(p_out &ImVec2, label &i8, has_close_button_or_unsaved_marker bool)

@[c: 'igTabItemCalcSize_WindowPtr']
pub fn tab_item_calc_size_window_ptr(p_out &ImVec2, window &Window)

@[c: 'igTabItemBackground']
pub fn tab_item_background(draw_list &ImDrawList, bb ImRect, flags TabItemFlags, col ImU32)

@[c: 'igTabItemLabelAndCloseButton']
pub fn tab_item_label_and_close_button(draw_list &ImDrawList, bb ImRect, flags TabItemFlags, frame_padding ImVec2, label &i8, tab_id ID, close_button_id ID, is_contents_visible bool, out_just_closed &bool, out_text_clipped &bool)

@[c: 'igRenderText']
pub fn render_text(pos ImVec2, text &i8, text_end &i8, hide_text_after_hash bool)

@[c: 'igRenderTextWrapped']
pub fn render_text_wrapped(pos ImVec2, text &i8, text_end &i8, wrap_width f32)

@[c: 'igRenderTextClipped']
pub fn render_text_clipped(pos_min ImVec2, pos_max ImVec2, text &i8, text_end &i8, text_size_if_known &ImVec2, align ImVec2, clip_rect &ImRect)

@[c: 'igRenderTextClippedEx']
pub fn render_text_clipped_ex(draw_list &ImDrawList, pos_min ImVec2, pos_max ImVec2, text &i8, text_end &i8, text_size_if_known &ImVec2, align ImVec2, clip_rect &ImRect)

@[c: 'igRenderTextEllipsis']
pub fn render_text_ellipsis(draw_list &ImDrawList, pos_min ImVec2, pos_max ImVec2, clip_max_x f32, ellipsis_max_x f32, text &i8, text_end &i8, text_size_if_known &ImVec2)

@[c: 'igRenderFrame']
pub fn render_frame(p_min ImVec2, p_max ImVec2, fill_col ImU32, borders bool, rounding f32)

@[c: 'igRenderFrameBorder']
pub fn render_frame_border(p_min ImVec2, p_max ImVec2, rounding f32)

@[c: 'igRenderColorRectWithAlphaCheckerboard']
pub fn render_color_rect_with_alpha_checkerboard(draw_list &ImDrawList, p_min ImVec2, p_max ImVec2, fill_col ImU32, grid_step f32, grid_off ImVec2, rounding f32, flags ImDrawFlags)

@[c: 'igRenderNavCursor']
pub fn render_nav_cursor(bb ImRect, id ID, flags NavRenderCursorFlags)

@[c: 'igFindRenderedTextEnd']
pub fn find_rendered_text_end(text &i8, text_end &i8) &i8

@[c: 'igRenderMouseCursor']
pub fn render_mouse_cursor(pos ImVec2, scale f32, mouse_cursor MouseCursor, col_fill ImU32, col_border ImU32, col_shadow ImU32)

@[c: 'igRenderArrow']
pub fn render_arrow(draw_list &ImDrawList, pos ImVec2, col ImU32, dir Dir, scale f32)

@[c: 'igRenderBullet']
pub fn render_bullet(draw_list &ImDrawList, pos ImVec2, col ImU32)

@[c: 'igRenderCheckMark']
pub fn render_check_mark(draw_list &ImDrawList, pos ImVec2, col ImU32, sz f32)

@[c: 'igRenderArrowPointingAt']
pub fn render_arrow_pointing_at(draw_list &ImDrawList, pos ImVec2, half_sz ImVec2, direction Dir, col ImU32)

@[c: 'igRenderArrowDockMenu']
pub fn render_arrow_dock_menu(draw_list &ImDrawList, p_min ImVec2, sz f32, col ImU32)

@[c: 'igRenderRectFilledRangeH']
pub fn render_rect_filled_range_h(draw_list &ImDrawList, rect ImRect, col ImU32, x_start_norm f32, x_end_norm f32, rounding f32)

@[c: 'igRenderRectFilledWithHole']
pub fn render_rect_filled_with_hole(draw_list &ImDrawList, outer ImRect, inner ImRect, col ImU32, rounding f32)

@[c: 'igCalcRoundingFlagsForRectInRect']
pub fn calc_rounding_flags_for_rect_in_rect(r_in ImRect, r_outer ImRect, threshold f32) ImDrawFlags

@[c: 'igTextEx']
pub fn text_ex(text &i8, text_end &i8, flags TextFlags)

@[c: 'igButtonEx']
pub fn button_ex(label &i8, size_arg ImVec2, flags ButtonFlags) bool

@[c: 'igArrowButtonEx']
pub fn arrow_button_ex(str_id &i8, dir Dir, size_arg ImVec2, flags ButtonFlags) bool

@[c: 'igImageButtonEx']
pub fn image_button_ex(id ID, user_texture_id ImTextureID, image_size ImVec2, uv0 ImVec2, uv1 ImVec2, bg_col ImVec4, tint_col ImVec4, flags ButtonFlags) bool

@[c: 'igSeparatorEx']
pub fn separator_ex(flags SeparatorFlags, thickness f32)

@[c: 'igSeparatorTextEx']
pub fn separator_text_ex(id ID, label &i8, label_end &i8, extra_width f32)

@[c: 'igCheckboxFlags_S64Ptr']
pub fn checkbox_flags_s64_ptr(label &i8, flags &ImS64, flags_value ImS64) bool

@[c: 'igCheckboxFlags_U64Ptr']
pub fn checkbox_flags_u64_ptr(label &i8, flags &ImU64, flags_value ImU64) bool

@[c: 'igCloseButton']
pub fn close_button(id ID, pos ImVec2) bool

@[c: 'igCollapseButton']
pub fn collapse_button(id ID, pos ImVec2, dock_node &DockNode) bool

@[c: 'igScrollbar']
pub fn scrollbar(axis Axis)

@[c: 'igScrollbarEx']
pub fn scrollbar_ex(bb ImRect, id ID, axis Axis, p_scroll_v &ImS64, avail_v ImS64, contents_v ImS64, draw_rounding_flags ImDrawFlags) bool

@[c: 'igGetWindowScrollbarRect']
pub fn get_window_scrollbar_rect(p_out &ImRect, window &Window, axis Axis)

@[c: 'igGetWindowScrollbarID']
pub fn get_window_scrollbar_id(window &Window, axis Axis) ID

@[c: 'igGetWindowResizeCornerID']
pub fn get_window_resize_corner_id(window &Window, n int) ID

@[c: 'igGetWindowResizeBorderID']
pub fn get_window_resize_border_id(window &Window, dir Dir) ID

@[c: 'igButtonBehavior']
pub fn button_behavior(bb ImRect, id ID, out_hovered &bool, out_held &bool, flags ButtonFlags) bool

@[c: 'igDragBehavior']
pub fn drag_behavior(id ID, data_type DataType, p_v voidptr, v_speed f32, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags) bool

@[c: 'igSliderBehavior']
pub fn slider_behavior(bb ImRect, id ID, data_type DataType, p_v voidptr, p_min voidptr, p_max voidptr, format &i8, flags SliderFlags, out_grab_bb &ImRect) bool

@[c: 'igSplitterBehavior']
pub fn splitter_behavior(bb ImRect, id ID, axis Axis, size1 &f32, size2 &f32, min_size1 f32, min_size2 f32, hover_extend f32, hover_visibility_delay f32, bg_col ImU32) bool

@[c: 'igTreeNodeBehavior']
pub fn tree_node_behavior(id ID, flags TreeNodeFlags, label &i8, label_end &i8) bool

@[c: 'igTreePushOverrideID']
pub fn tree_push_override_id(id ID)

@[c: 'igTreeNodeGetOpen']
pub fn tree_node_get_open(storage_id ID) bool

@[c: 'igTreeNodeSetOpen']
pub fn tree_node_set_open(storage_id ID, open bool)

@[c: 'igTreeNodeUpdateNextOpen']
pub fn tree_node_update_next_open(storage_id ID, flags TreeNodeFlags) bool

@[c: 'igDataTypeGetInfo']
pub fn data_type_get_info(data_type DataType) &DataTypeInfo

@[c: 'igDataTypeFormatString']
pub fn data_type_format_string(buf &i8, buf_size int, data_type DataType, p_data voidptr, format &i8) int

@[c: 'igDataTypeApplyOp']
pub fn data_type_apply_op(data_type DataType, op int, output voidptr, arg_1 voidptr, arg_2 voidptr)

@[c: 'igDataTypeApplyFromText']
pub fn data_type_apply_from_text(buf &i8, data_type DataType, p_data voidptr, format &i8, p_data_when_empty voidptr) bool

@[c: 'igDataTypeCompare']
pub fn data_type_compare(data_type DataType, arg_1 voidptr, arg_2 voidptr) int

@[c: 'igDataTypeClamp']
pub fn data_type_clamp(data_type DataType, p_data voidptr, p_min voidptr, p_max voidptr) bool

@[c: 'igDataTypeIsZero']
pub fn data_type_is_zero(data_type DataType, p_data voidptr) bool

@[c: 'igInputTextEx']
pub fn input_text_ex(label &i8, hint &i8, buf &i8, buf_size int, size_arg ImVec2, flags InputTextFlags, callback InputTextCallback, user_data voidptr) bool

@[c: 'igInputTextDeactivateHook']
pub fn input_text_deactivate_hook(id ID)

@[c: 'igTempInputText']
pub fn temp_input_text(bb ImRect, id ID, label &i8, buf &i8, buf_size int, flags InputTextFlags) bool

@[c: 'igTempInputScalar']
pub fn temp_input_scalar(bb ImRect, id ID, label &i8, data_type DataType, p_data voidptr, format &i8, p_clamp_min voidptr, p_clamp_max voidptr) bool

@[c: 'igTempInputIsActive']
pub fn temp_input_is_active(id ID) bool

@[c: 'igGetInputTextState']
pub fn get_input_text_state(id ID) &InputTextState

@[c: 'igSetNextItemRefVal']
pub fn set_next_item_ref_val(data_type DataType, p_data voidptr)

@[c: 'igIsItemActiveAsInputText']
pub fn is_item_active_as_input_text() bool

@[c: 'igColorTooltip']
pub fn color_tooltip(text &i8, col &f32, flags ColorEditFlags)

@[c: 'igColorEditOptionsPopup']
pub fn color_edit_options_popup(col &f32, flags ColorEditFlags)

@[c: 'igColorPickerOptionsPopup']
pub fn color_picker_options_popup(ref_col &f32, flags ColorEditFlags)

@[c: 'igPlotEx']
pub fn plot_ex(plot_type PlotType, label &i8, values_getter fn (voidptr, int) f32, data voidptr, values_count int, values_offset int, overlay_text &i8, scale_min f32, scale_max f32, size_arg ImVec2) int

@[c: 'igShadeVertsLinearColorGradientKeepAlpha']
pub fn shade_verts_linear_color_gradient_keep_alpha(draw_list &ImDrawList, vert_start_idx int, vert_end_idx int, gradient_p0 ImVec2, gradient_p1 ImVec2, col0 ImU32, col1 ImU32)

@[c: 'igShadeVertsLinearUV']
pub fn shade_verts_linear_uv(draw_list &ImDrawList, vert_start_idx int, vert_end_idx int, a ImVec2, b ImVec2, uv_a ImVec2, uv_b ImVec2, clamp bool)

@[c: 'igShadeVertsTransformPos']
pub fn shade_verts_transform_pos(draw_list &ImDrawList, vert_start_idx int, vert_end_idx int, pivot_in ImVec2, cos_a f32, sin_a f32, pivot_out ImVec2)

@[c: 'igGcCompactTransientMiscBuffers']
pub fn gc_compact_transient_misc_buffers()

@[c: 'igGcCompactTransientWindowBuffers']
pub fn gc_compact_transient_window_buffers(window &Window)

@[c: 'igGcAwakeTransientWindowBuffers']
pub fn gc_awake_transient_window_buffers(window &Window)

@[c: 'igErrorLog']
pub fn error_log(msg &i8) bool

@[c: 'igErrorRecoveryStoreState']
pub fn error_recovery_store_state(state_out &ErrorRecoveryState)

@[c: 'igErrorRecoveryTryToRecoverState']
pub fn error_recovery_try_to_recover_state(state_in &ErrorRecoveryState)

@[c: 'igErrorRecoveryTryToRecoverWindowState']
pub fn error_recovery_try_to_recover_window_state(state_in &ErrorRecoveryState)

@[c: 'igErrorCheckUsingSetCursorPosToExtendParentBoundaries']
pub fn error_check_using_set_cursor_pos_to_extend_parent_boundaries()

@[c: 'igErrorCheckEndFrameFinalizeErrorTooltip']
pub fn error_check_end_frame_finalize_error_tooltip()

@[c: 'igBeginErrorTooltip']
pub fn begin_error_tooltip() bool

@[c: 'igEndErrorTooltip']
pub fn end_error_tooltip()

@[c: 'igDebugAllocHook']
pub fn debug_alloc_hook(info &DebugAllocInfo, frame_count int, ptr voidptr, size usize)

@[c: 'igDebugDrawCursorPos']
pub fn debug_draw_cursor_pos(col ImU32)

@[c: 'igDebugDrawLineExtents']
pub fn debug_draw_line_extents(col ImU32)

@[c: 'igDebugDrawItemRect']
pub fn debug_draw_item_rect(col ImU32)

@[c: 'igDebugTextUnformattedWithLocateItem']
pub fn debug_text_unformatted_with_locate_item(line_begin &i8, line_end &i8)

@[c: 'igDebugLocateItem']
pub fn debug_locate_item(target_id ID)

@[c: 'igDebugLocateItemOnHover']
pub fn debug_locate_item_on_hover(target_id ID)

@[c: 'igDebugLocateItemResolveWithLastItem']
pub fn debug_locate_item_resolve_with_last_item()

@[c: 'igDebugBreakClearData']
pub fn debug_break_clear_data()

@[c: 'igDebugBreakButton']
pub fn debug_break_button(label &i8, description_of_location &i8) bool

@[c: 'igDebugBreakButtonTooltip']
pub fn debug_break_button_tooltip(keyboard_only bool, description_of_location &i8)

@[c: 'igShowFontAtlas']
pub fn show_font_atlas(atlas &ImFontAtlas)

@[c: 'igDebugHookIdInfo']
pub fn debug_hook_id_info(id ID, data_type DataType, data_id voidptr, data_id_end voidptr)

@[c: 'igDebugNodeColumns']
pub fn debug_node_columns(columns &OldColumns)

@[c: 'igDebugNodeDockNode']
pub fn debug_node_dock_node(node &DockNode, label &i8)

@[c: 'igDebugNodeDrawList']
pub fn debug_node_draw_list(window &Window, viewport &ViewportP, draw_list &ImDrawList, label &i8)

@[c: 'igDebugNodeDrawCmdShowMeshAndBoundingBox']
pub fn debug_node_draw_cmd_show_mesh_and_bounding_box(out_draw_list &ImDrawList, draw_list &ImDrawList, draw_cmd &ImDrawCmd, show_mesh bool, show_aabb bool)

@[c: 'igDebugNodeFont']
pub fn debug_node_font(font &ImFont)

@[c: 'igDebugNodeFontGlyph']
pub fn debug_node_font_glyph(font &ImFont, glyph &ImFontGlyph)

@[c: 'igDebugNodeStorage']
pub fn debug_node_storage(storage &Storage, label &i8)

@[c: 'igDebugNodeTabBar']
pub fn debug_node_tab_bar(tab_bar &TabBar, label &i8)

@[c: 'igDebugNodeTable']
pub fn debug_node_table(table &Table)

@[c: 'igDebugNodeTableSettings']
pub fn debug_node_table_settings(settings &TableSettings)

@[c: 'igDebugNodeInputTextState']
pub fn debug_node_input_text_state(state &InputTextState)

@[c: 'igDebugNodeTypingSelectState']
pub fn debug_node_typing_select_state(state &TypingSelectState)

@[c: 'igDebugNodeMultiSelectState']
pub fn debug_node_multi_select_state(state &MultiSelectState)

@[c: 'igDebugNodeWindow']
pub fn debug_node_window(window &Window, label &i8)

@[c: 'igDebugNodeWindowSettings']
pub fn debug_node_window_settings(settings &WindowSettings)

@[c: 'igDebugNodeWindowsList']
pub fn debug_node_windows_list(windows &ImVector_WindowPtr, label &i8)

@[c: 'igDebugNodeWindowsListByBeginStackParent']
pub fn debug_node_windows_list_by_begin_stack_parent(windows &&Window, windows_size int, parent_in_begin_stack &Window)

@[c: 'igDebugNodeViewport']
pub fn debug_node_viewport(viewport &ViewportP)

@[c: 'igDebugNodePlatformMonitor']
pub fn debug_node_platform_monitor(monitor &PlatformMonitor, label &i8, idx int)

@[c: 'igDebugRenderKeyboardPreview']
pub fn debug_render_keyboard_preview(draw_list &ImDrawList)

@[c: 'igDebugRenderViewportThumbnail']
pub fn debug_render_viewport_thumbnail(draw_list &ImDrawList, viewport &ViewportP, bb ImRect)

@[c: 'igImFontAtlasGetBuilderForStbTruetype']
pub fn im_font_atlas_get_builder_for_stb_truetype() &ImFontBuilderIO

@[c: 'igImFontAtlasUpdateSourcesPointers']
pub fn im_font_atlas_update_sources_pointers(atlas &ImFontAtlas)

@[c: 'igImFontAtlasBuildInit']
pub fn im_font_atlas_build_init(atlas &ImFontAtlas)

@[c: 'igImFontAtlasBuildSetupFont']
pub fn im_font_atlas_build_setup_font(atlas &ImFontAtlas, font &ImFont, src &ImFontConfig, ascent f32, descent f32)

@[c: 'igImFontAtlasBuildPackCustomRects']
pub fn im_font_atlas_build_pack_custom_rects(atlas &ImFontAtlas, stbrp_context_opaque voidptr)

@[c: 'igImFontAtlasBuildFinish']
pub fn im_font_atlas_build_finish(atlas &ImFontAtlas)

@[c: 'igImFontAtlasBuildRender8bppRectFromString']
pub fn im_font_atlas_build_render8bpp_rect_from_string(atlas &ImFontAtlas, x int, y int, w int, h int, in_str &i8, in_marker_char i8, in_marker_pixel_value u8)

@[c: 'igImFontAtlasBuildRender32bppRectFromString']
pub fn im_font_atlas_build_render32bpp_rect_from_string(atlas &ImFontAtlas, x int, y int, w int, h int, in_str &i8, in_marker_char i8, in_marker_pixel_value u32)

@[c: 'igImFontAtlasBuildMultiplyCalcLookupTable']
pub fn im_font_atlas_build_multiply_calc_lookup_table(out_table &u8, in_multiply_factor f32)

@[c: 'igImFontAtlasBuildMultiplyRectAlpha8']
pub fn im_font_atlas_build_multiply_rect_alpha8(table &u8, pixels &u8, x int, y int, w int, h int, stride int)

@[c: 'igImFontAtlasBuildGetOversampleFactors']
pub fn im_font_atlas_build_get_oversample_factors(src &ImFontConfig, out_oversample_h &int, out_oversample_v &int)

@[c: 'igImFontAtlasGetMouseCursorTexData']
pub fn im_font_atlas_get_mouse_cursor_tex_data(atlas &ImFontAtlas, cursor_type MouseCursor, out_offset &ImVec2, out_size &ImVec2, out_uv_border &ImVec2, out_uv_fill &ImVec2) bool

/////////////////////////hand written functions
// no LogTextV
@[c: 'igLogText']
@[c2v_variadic]
pub fn log_text(fmt ...&i8)

// no appendfV
@[c: 'TextBuffer_appendf']
@[c2v_variadic]
pub fn text_buffer_appendf(self &TextBuffer, fmt ...&i8)

// for getting FLT_MAX in bindings
@[c: 'igGET_FLT_MAX']
pub fn get_flt_max() f32

// for getting FLT_MIN in bindings
@[c: 'igGET_FLT_MIN']
pub fn get_flt_min() f32

@[c: 'ImVector_ImWchar_create']
pub fn im_vector_im_wchar_create() &ImVector_ImWchar

@[c: 'ImVector_ImWchar_destroy']
pub fn im_vector_im_wchar_destroy(self &ImVector_ImWchar)

@[c: 'ImVector_ImWchar_Init']
pub fn im_vector_im_wchar_init(p &ImVector_ImWchar)

@[c: 'ImVector_ImWchar_UnInit']
pub fn im_vector_im_wchar_un_init(p &ImVector_ImWchar)

@[c: 'PlatformIO_Set_Platform_GetWindowPos']
pub fn platform_io_set_platform_get_window_pos(platform_io &PlatformIO, user_callback fn (&Viewport, ImVec2))

@[c: 'PlatformIO_Set_Platform_GetWindowSize']
pub fn platform_io_set_platform_get_window_size(platform_io &PlatformIO, user_callback fn (&Viewport, ImVec2))

// CIMGUI_INCLUDED
